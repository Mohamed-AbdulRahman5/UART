
module tx_D_bits9_sb_tick16 ( clk, reset_n, data_in, tx_start, s_tick, tx, 
        tx_done, parity_bit );
  input [7:0] data_in;
  input clk, reset_n, tx_start, s_tick;
  output tx, tx_done, parity_bit;
  wire   n2, n4, n5, n9, n10, n11, n13, n16, n19, n20, n21, n23, n25, n27, n29,
         n31, n34, n36, n37, n38, n39, n40, n41, n42, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n66, n67, n71, n74, n81, n82, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188;

  XOR2_X1 U58 ( .A(n60), .B(n61), .Z(n46) );
  DFF_X1 tx_reg ( .D(n82), .CK(clk), .Q(tx), .QN(n188) );
  DFFR_X1 state_reg_reg_0_ ( .D(n110), .CK(clk), .RN(reset_n), .Q(n176), .QN(
        n96) );
  DFFR_X1 state_reg_reg_1_ ( .D(n113), .CK(clk), .RN(reset_n), .Q(n179), .QN(
        n95) );
  DFFR_X1 s_reg_reg_2_ ( .D(n112), .CK(clk), .RN(reset_n), .QN(n97) );
  DFFR_X1 n_reg_reg_2_ ( .D(n107), .CK(clk), .RN(reset_n), .QN(n91) );
  DFFR_X1 n_reg_reg_1_ ( .D(n108), .CK(clk), .RN(reset_n), .QN(n92) );
  DFFR_X1 n_reg_reg_0_ ( .D(n109), .CK(clk), .RN(reset_n), .QN(n93) );
  DFFR_X1 b_reg_reg_7_ ( .D(n163), .CK(clk), .RN(reset_n), .Q(n180) );
  DFFR_X1 b_reg_reg_6_ ( .D(n99), .CK(clk), .RN(reset_n), .Q(n181), .QN(n84)
         );
  DFFR_X1 b_reg_reg_5_ ( .D(n100), .CK(clk), .RN(reset_n), .Q(n182), .QN(n85)
         );
  DFFR_X1 b_reg_reg_4_ ( .D(n101), .CK(clk), .RN(reset_n), .Q(n183), .QN(n86)
         );
  DFFR_X1 b_reg_reg_3_ ( .D(n102), .CK(clk), .RN(reset_n), .Q(n184), .QN(n87)
         );
  DFFR_X1 b_reg_reg_2_ ( .D(n103), .CK(clk), .RN(reset_n), .Q(n185), .QN(n88)
         );
  DFFR_X1 b_reg_reg_1_ ( .D(n104), .CK(clk), .RN(reset_n), .Q(n186), .QN(n89)
         );
  DFFR_X1 b_reg_reg_0_ ( .D(n105), .CK(clk), .RN(reset_n), .QN(n90) );
  DFFR_X1 s_reg_reg_3_ ( .D(n114), .CK(clk), .RN(reset_n), .QN(n172) );
  DFFR_X1 s_reg_reg_1_ ( .D(n111), .CK(clk), .RN(reset_n), .QN(n187) );
  DFFR_X1 s_reg_reg_0_ ( .D(n115), .CK(clk), .RN(reset_n), .QN(n171) );
  DFFR_X1 n_reg_reg_3_ ( .D(n106), .CK(clk), .RN(reset_n), .Q(n81), .QN(n173)
         );
  DFFR_X1 parity_bit_reg ( .D(n98), .CK(clk), .RN(reset_n), .Q(parity_bit) );
  NAND2_X1 U3 ( .A1(n169), .A2(n165), .ZN(n45) );
  INV_X1 U4 ( .A(n71), .ZN(n168) );
  INV_X1 U5 ( .A(n49), .ZN(n169) );
  AND2_X1 U6 ( .A1(n178), .A2(n34), .ZN(n10) );
  INV_X1 U7 ( .A(n11), .ZN(n164) );
  AND2_X1 U8 ( .A1(n169), .A2(n34), .ZN(n20) );
  NOR2_X1 U9 ( .A1(n177), .A2(n54), .ZN(n53) );
  NAND2_X1 U10 ( .A1(n57), .A2(n71), .ZN(n58) );
  INV_X1 U11 ( .A(s_tick), .ZN(n166) );
  NAND2_X1 U12 ( .A1(n177), .A2(n166), .ZN(n39) );
  INV_X1 U13 ( .A(n37), .ZN(n165) );
  NAND2_X1 U14 ( .A1(n16), .A2(n177), .ZN(n49) );
  NOR2_X1 U15 ( .A1(n170), .A2(n174), .ZN(n16) );
  OAI21_X1 U16 ( .B1(n177), .B2(n175), .A(n170), .ZN(n51) );
  NAND2_X1 U17 ( .A1(n51), .A2(n41), .ZN(n71) );
  OR2_X1 U18 ( .A1(n41), .A2(n170), .ZN(n13) );
  NAND4_X1 U19 ( .A1(n39), .A2(n40), .A3(n52), .A4(n41), .ZN(n37) );
  NAND2_X1 U20 ( .A1(n62), .A2(n74), .ZN(n57) );
  NAND3_X1 U21 ( .A1(n13), .A2(n52), .A3(s_tick), .ZN(n74) );
  OAI21_X1 U22 ( .B1(n16), .B2(n36), .A(n34), .ZN(n11) );
  OAI22_X1 U23 ( .A1(n171), .A2(n57), .B1(n48), .B2(n58), .ZN(n115) );
  AND2_X1 U24 ( .A1(n62), .A2(n63), .ZN(n54) );
  NAND3_X1 U25 ( .A1(n64), .A2(n52), .A3(s_tick), .ZN(n63) );
  OAI22_X1 U26 ( .A1(n187), .A2(n57), .B1(n47), .B2(n58), .ZN(n111) );
  OAI22_X1 U27 ( .A1(n172), .A2(n57), .B1(n44), .B2(n58), .ZN(n114) );
  OAI22_X1 U28 ( .A1(n42), .A2(n173), .B1(n44), .B2(n45), .ZN(n106) );
  NAND2_X1 U29 ( .A1(n37), .A2(n38), .ZN(n34) );
  NAND4_X1 U30 ( .A1(tx_start), .A2(n39), .A3(n40), .A4(n41), .ZN(n38) );
  AND2_X1 U31 ( .A1(n50), .A2(n51), .ZN(n42) );
  OAI21_X1 U32 ( .B1(n166), .B2(n40), .A(n37), .ZN(n50) );
  NOR2_X1 U33 ( .A1(n13), .A2(n166), .ZN(tx_done) );
  INV_X1 U34 ( .A(n9), .ZN(n163) );
  AOI22_X1 U35 ( .A1(data_in[7]), .A2(n10), .B1(n11), .B2(n180), .ZN(n9) );
  INV_X1 U36 ( .A(n36), .ZN(n177) );
  OAI21_X1 U37 ( .B1(n59), .B2(n48), .A(n60), .ZN(n47) );
  XNOR2_X1 U38 ( .A(n66), .B(n67), .ZN(n44) );
  OAI22_X1 U39 ( .A1(n173), .A2(n49), .B1(n168), .B2(n172), .ZN(n66) );
  NOR2_X1 U40 ( .A1(n167), .A2(n60), .ZN(n67) );
  INV_X1 U41 ( .A(n61), .ZN(n167) );
  NAND2_X1 U42 ( .A1(n48), .A2(n59), .ZN(n60) );
  NAND2_X1 U43 ( .A1(n176), .A2(n179), .ZN(n41) );
  INV_X1 U44 ( .A(n64), .ZN(n170) );
  INV_X1 U45 ( .A(n5), .ZN(n174) );
  INV_X1 U46 ( .A(n40), .ZN(n175) );
  INV_X1 U47 ( .A(n52), .ZN(n178) );
  OAI21_X1 U48 ( .B1(n90), .B2(n164), .A(n31), .ZN(n105) );
  AOI22_X1 U49 ( .A1(data_in[0]), .A2(n10), .B1(n20), .B2(n186), .ZN(n31) );
  OAI21_X1 U50 ( .B1(n89), .B2(n164), .A(n29), .ZN(n104) );
  AOI22_X1 U51 ( .A1(data_in[1]), .A2(n10), .B1(n20), .B2(n185), .ZN(n29) );
  OAI21_X1 U52 ( .B1(n88), .B2(n164), .A(n27), .ZN(n103) );
  AOI22_X1 U53 ( .A1(data_in[2]), .A2(n10), .B1(n20), .B2(n184), .ZN(n27) );
  OAI21_X1 U54 ( .B1(n87), .B2(n164), .A(n25), .ZN(n102) );
  AOI22_X1 U55 ( .A1(data_in[3]), .A2(n10), .B1(n20), .B2(n183), .ZN(n25) );
  OAI21_X1 U56 ( .B1(n86), .B2(n164), .A(n23), .ZN(n101) );
  AOI22_X1 U57 ( .A1(data_in[4]), .A2(n10), .B1(n20), .B2(n182), .ZN(n23) );
  OAI21_X1 U59 ( .B1(n85), .B2(n164), .A(n21), .ZN(n100) );
  AOI22_X1 U60 ( .A1(data_in[5]), .A2(n10), .B1(n20), .B2(n181), .ZN(n21) );
  OAI21_X1 U61 ( .B1(n84), .B2(n164), .A(n19), .ZN(n99) );
  AOI22_X1 U62 ( .A1(data_in[6]), .A2(n10), .B1(n20), .B2(n180), .ZN(n19) );
  OAI22_X1 U63 ( .A1(n54), .A2(n40), .B1(n95), .B2(n53), .ZN(n113) );
  OAI22_X1 U64 ( .A1(n93), .A2(n42), .B1(n45), .B2(n48), .ZN(n109) );
  OAI22_X1 U65 ( .A1(n97), .A2(n57), .B1(n46), .B2(n58), .ZN(n112) );
  OAI22_X1 U66 ( .A1(n91), .A2(n42), .B1(n45), .B2(n46), .ZN(n107) );
  OAI22_X1 U67 ( .A1(n96), .A2(n53), .B1(n54), .B2(n55), .ZN(n110) );
  AOI21_X1 U68 ( .B1(n174), .B2(n177), .A(n178), .ZN(n55) );
  OAI22_X1 U69 ( .A1(n92), .A2(n42), .B1(n45), .B2(n47), .ZN(n108) );
  XNOR2_X1 U70 ( .A(parity_bit), .B(n162), .ZN(n98) );
  NAND3_X1 U71 ( .A1(n16), .A2(n165), .A3(tx), .ZN(n162) );
  OAI21_X1 U72 ( .B1(reset_n), .B2(n188), .A(n2), .ZN(n82) );
  OAI221_X1 U73 ( .B1(n174), .B2(n4), .C1(n5), .C2(parity_bit), .A(reset_n), 
        .ZN(n2) );
  AOI21_X1 U74 ( .B1(n90), .B2(n177), .A(n175), .ZN(n4) );
  NOR4_X1 U75 ( .A1(n171), .A2(n172), .A3(n187), .A4(n97), .ZN(n64) );
  OAI22_X1 U76 ( .A1(n93), .A2(n49), .B1(n168), .B2(n171), .ZN(n48) );
  NAND2_X1 U77 ( .A1(n95), .A2(n176), .ZN(n40) );
  OAI22_X1 U78 ( .A1(n92), .A2(n49), .B1(n168), .B2(n187), .ZN(n59) );
  OAI22_X1 U79 ( .A1(n91), .A2(n49), .B1(n168), .B2(n97), .ZN(n61) );
  NAND4_X1 U80 ( .A1(n81), .A2(n91), .A3(n92), .A4(n93), .ZN(n5) );
  NAND3_X1 U81 ( .A1(n95), .A2(n40), .A3(tx_start), .ZN(n62) );
  NAND2_X1 U82 ( .A1(n96), .A2(n179), .ZN(n36) );
  NAND2_X1 U83 ( .A1(n95), .A2(n96), .ZN(n52) );
endmodule


module dual_gray_counter_addr_size8_1_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[8]), .B(A[8]), .Z(SUM[8]) );
endmodule


module dual_gray_counter_addr_size8_1 ( clk, gray_count_st, gray_count_nd, 
        reset_n, en );
  output [8:0] gray_count_st;
  output [7:0] gray_count_nd;
  input clk, reset_n, en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [7:0] Q_reg;
  wire   [8:0] Q_next;
  assign gray_count_nd[6] = gray_count_st[6];
  assign gray_count_nd[5] = gray_count_st[5];
  assign gray_count_nd[4] = gray_count_st[4];
  assign gray_count_nd[3] = gray_count_st[3];
  assign gray_count_nd[1] = gray_count_st[1];
  assign gray_count_nd[0] = gray_count_st[0];
  assign gray_count_nd[2] = gray_count_st[2];

  XOR2_X1 U22 ( .A(n12), .B(n13), .Z(gray_count_st[5]) );
  XOR2_X1 U23 ( .A(n13), .B(n14), .Z(gray_count_st[4]) );
  XOR2_X1 U24 ( .A(n14), .B(n15), .Z(gray_count_st[3]) );
  XOR2_X1 U26 ( .A(n16), .B(n17), .Z(gray_count_st[1]) );
  XOR2_X1 U29 ( .A(n11), .B(n10), .Z(gray_count_st[7]) );
  dual_gray_counter_addr_size8_1_DW01_inc_0 add_48 ( .A({gray_count_st[8], 
        Q_reg}), .SUM(Q_next) );
  DFFR_X1 Q_reg_reg_8_ ( .D(n19), .CK(clk), .RN(reset_n), .Q(gray_count_st[8]), 
        .QN(n10) );
  DFFR_X1 Q_reg_reg_7_ ( .D(n20), .CK(clk), .RN(reset_n), .Q(Q_reg[7]), .QN(
        n11) );
  DFFR_X1 Q_reg_reg_6_ ( .D(n21), .CK(clk), .RN(reset_n), .Q(Q_reg[6]), .QN(
        n12) );
  DFFR_X1 Q_reg_reg_5_ ( .D(n22), .CK(clk), .RN(reset_n), .Q(Q_reg[5]), .QN(
        n13) );
  DFFR_X1 Q_reg_reg_4_ ( .D(n23), .CK(clk), .RN(reset_n), .Q(Q_reg[4]), .QN(
        n14) );
  DFFR_X1 Q_reg_reg_3_ ( .D(n24), .CK(clk), .RN(reset_n), .Q(Q_reg[3]), .QN(
        n15) );
  DFFR_X1 Q_reg_reg_2_ ( .D(n25), .CK(clk), .RN(reset_n), .Q(Q_reg[2]), .QN(
        n16) );
  DFFR_X1 Q_reg_reg_1_ ( .D(n26), .CK(clk), .RN(reset_n), .Q(Q_reg[1]), .QN(
        n17) );
  DFFR_X1 Q_reg_reg_0_ ( .D(n27), .CK(clk), .RN(reset_n), .Q(Q_reg[0]), .QN(
        n18) );
  XNOR2_X1 U3 ( .A(Q_reg[1]), .B(n18), .ZN(gray_count_st[0]) );
  XNOR2_X1 U4 ( .A(Q_reg[3]), .B(n16), .ZN(gray_count_st[2]) );
  XOR2_X2 U5 ( .A(n11), .B(n12), .Z(gray_count_st[6]) );
  OAI21_X1 U6 ( .B1(n10), .B2(en), .A(n1), .ZN(n19) );
  NAND2_X1 U7 ( .A1(en), .A2(Q_next[8]), .ZN(n1) );
  OAI21_X1 U8 ( .B1(n11), .B2(en), .A(n2), .ZN(n20) );
  NAND2_X1 U9 ( .A1(Q_next[7]), .A2(en), .ZN(n2) );
  OAI21_X1 U10 ( .B1(n12), .B2(en), .A(n3), .ZN(n21) );
  NAND2_X1 U11 ( .A1(Q_next[6]), .A2(en), .ZN(n3) );
  OAI21_X1 U12 ( .B1(n13), .B2(en), .A(n4), .ZN(n22) );
  NAND2_X1 U13 ( .A1(Q_next[5]), .A2(en), .ZN(n4) );
  OAI21_X1 U14 ( .B1(n14), .B2(en), .A(n5), .ZN(n23) );
  NAND2_X1 U15 ( .A1(Q_next[4]), .A2(en), .ZN(n5) );
  OAI21_X1 U16 ( .B1(n15), .B2(en), .A(n6), .ZN(n24) );
  NAND2_X1 U17 ( .A1(Q_next[3]), .A2(en), .ZN(n6) );
  OAI21_X1 U18 ( .B1(n16), .B2(en), .A(n7), .ZN(n25) );
  NAND2_X1 U19 ( .A1(Q_next[2]), .A2(en), .ZN(n7) );
  OAI21_X1 U20 ( .B1(n17), .B2(en), .A(n8), .ZN(n26) );
  NAND2_X1 U21 ( .A1(Q_next[1]), .A2(en), .ZN(n8) );
  OAI21_X1 U25 ( .B1(n18), .B2(en), .A(n9), .ZN(n27) );
  NAND2_X1 U27 ( .A1(Q_next[0]), .A2(en), .ZN(n9) );
  XNOR2_X1 U28 ( .A(n10), .B(gray_count_st[7]), .ZN(gray_count_nd[7]) );
endmodule


module dual_gray_counter_addr_size8_3_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[8]), .B(A[8]), .Z(SUM[8]) );
endmodule


module dual_gray_counter_addr_size8_3 ( clk, gray_count_st, gray_count_nd, 
        reset_n, en );
  output [8:0] gray_count_st;
  output [7:0] gray_count_nd;
  input clk, reset_n, en;
  wire   n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55;
  wire   [7:0] Q_reg;
  wire   [8:0] Q_next;
  assign gray_count_nd[6] = gray_count_st[6];
  assign gray_count_nd[5] = gray_count_st[5];
  assign gray_count_nd[4] = gray_count_st[4];
  assign gray_count_nd[3] = gray_count_st[3];
  assign gray_count_nd[2] = gray_count_st[2];
  assign gray_count_nd[1] = gray_count_st[1];
  assign gray_count_nd[0] = gray_count_st[0];

  DFFR_X1 Q_reg_reg_0_ ( .D(n29), .CK(clk), .RN(reset_n), .Q(Q_reg[0]), .QN(
        n38) );
  DFFR_X1 Q_reg_reg_1_ ( .D(n30), .CK(clk), .RN(reset_n), .Q(Q_reg[1]), .QN(
        n39) );
  DFFR_X1 Q_reg_reg_2_ ( .D(n31), .CK(clk), .RN(reset_n), .Q(Q_reg[2]), .QN(
        n40) );
  DFFR_X1 Q_reg_reg_3_ ( .D(n32), .CK(clk), .RN(reset_n), .Q(Q_reg[3]), .QN(
        n41) );
  DFFR_X1 Q_reg_reg_4_ ( .D(n33), .CK(clk), .RN(reset_n), .Q(Q_reg[4]), .QN(
        n42) );
  DFFR_X1 Q_reg_reg_5_ ( .D(n34), .CK(clk), .RN(reset_n), .Q(Q_reg[5]), .QN(
        n43) );
  DFFR_X1 Q_reg_reg_6_ ( .D(n35), .CK(clk), .RN(reset_n), .Q(Q_reg[6]), .QN(
        n44) );
  DFFR_X1 Q_reg_reg_7_ ( .D(n36), .CK(clk), .RN(reset_n), .Q(Q_reg[7]), .QN(
        n45) );
  DFFR_X1 Q_reg_reg_8_ ( .D(n37), .CK(clk), .RN(reset_n), .Q(gray_count_st[8]), 
        .QN(n46) );
  XOR2_X1 U21 ( .A(n45), .B(n44), .Z(gray_count_st[6]) );
  XOR2_X1 U22 ( .A(n44), .B(n43), .Z(gray_count_st[5]) );
  XOR2_X1 U23 ( .A(n43), .B(n42), .Z(gray_count_st[4]) );
  XOR2_X1 U24 ( .A(n42), .B(n41), .Z(gray_count_st[3]) );
  XOR2_X1 U25 ( .A(n41), .B(n40), .Z(gray_count_st[2]) );
  XOR2_X1 U26 ( .A(n40), .B(n39), .Z(gray_count_st[1]) );
  XOR2_X1 U27 ( .A(n39), .B(n38), .Z(gray_count_st[0]) );
  XOR2_X1 U29 ( .A(n45), .B(n46), .Z(gray_count_st[7]) );
  dual_gray_counter_addr_size8_3_DW01_inc_0 add_48 ( .A({gray_count_st[8], 
        Q_reg}), .SUM(Q_next) );
  BUF_X1 U3 ( .A(en), .Z(n28) );
  OAI21_X1 U4 ( .B1(n44), .B2(en), .A(n53), .ZN(n35) );
  NAND2_X1 U5 ( .A1(Q_next[6]), .A2(n28), .ZN(n53) );
  OAI21_X1 U6 ( .B1(n43), .B2(en), .A(n52), .ZN(n34) );
  NAND2_X1 U7 ( .A1(Q_next[5]), .A2(n28), .ZN(n52) );
  OAI21_X1 U8 ( .B1(n42), .B2(en), .A(n51), .ZN(n33) );
  NAND2_X1 U9 ( .A1(Q_next[4]), .A2(n28), .ZN(n51) );
  OAI21_X1 U10 ( .B1(n41), .B2(en), .A(n50), .ZN(n32) );
  NAND2_X1 U11 ( .A1(Q_next[3]), .A2(n28), .ZN(n50) );
  OAI21_X1 U12 ( .B1(n40), .B2(n28), .A(n49), .ZN(n31) );
  NAND2_X1 U13 ( .A1(Q_next[2]), .A2(n28), .ZN(n49) );
  OAI21_X1 U14 ( .B1(n39), .B2(n28), .A(n48), .ZN(n30) );
  NAND2_X1 U15 ( .A1(Q_next[1]), .A2(n28), .ZN(n48) );
  OAI21_X1 U16 ( .B1(n45), .B2(en), .A(n54), .ZN(n36) );
  NAND2_X1 U17 ( .A1(Q_next[7]), .A2(n28), .ZN(n54) );
  OAI21_X1 U18 ( .B1(n46), .B2(n28), .A(n55), .ZN(n37) );
  NAND2_X1 U19 ( .A1(en), .A2(Q_next[8]), .ZN(n55) );
  OAI21_X1 U20 ( .B1(n38), .B2(n28), .A(n47), .ZN(n29) );
  NAND2_X1 U28 ( .A1(Q_next[0]), .A2(n28), .ZN(n47) );
  XNOR2_X1 U30 ( .A(n46), .B(gray_count_st[7]), .ZN(gray_count_nd[7]) );
endmodule


module fifo_control_unit_addr_size8_1 ( reset_n, w_clk, r_clk, rd, wr, addr_r, 
        addr_w, full, empty, we_enable, rd_enable );
  output [7:0] addr_r;
  output [7:0] addr_w;
  input reset_n, w_clk, r_clk, rd, wr;
  output full, empty, we_enable, rd_enable;
  wire   N4, n3, n40, n5, n1, n2, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n34;
  wire   [8:0] ptr_r;
  wire   [8:0] ptr_w;
  wire   [8:0] ptr_w_syn;
  wire   [8:0] ptr_w_syn_1;
  wire   [8:1] ptr_r_syn;
  wire   [8:0] ptr_r_syn_1;

  NOR2_X2 U4 ( .A1(empty), .A2(n34), .ZN(rd_enable) );
  XOR2_X1 U8 ( .A(ptr_w[8]), .B(ptr_r_syn[8]), .Z(n5) );
  XOR2_X1 U9 ( .A(ptr_w[7]), .B(ptr_r_syn[7]), .Z(n40) );
  dual_gray_counter_addr_size8_1 read_ptr ( .clk(r_clk), .gray_count_st(ptr_r), 
        .gray_count_nd(addr_r), .reset_n(reset_n), .en(rd_enable) );
  dual_gray_counter_addr_size8_3 write_ptr ( .clk(w_clk), .gray_count_st(ptr_w), .gray_count_nd(addr_w), .reset_n(reset_n), .en(we_enable) );
  DFFR_X1 ptr_w_syn_reg_8_ ( .D(ptr_w_syn_1[8]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[8]) );
  DFFR_X1 ptr_w_syn_reg_7_ ( .D(ptr_w_syn_1[7]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[7]) );
  DFFR_X1 ptr_w_syn_reg_6_ ( .D(ptr_w_syn_1[6]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[6]) );
  DFFR_X1 ptr_w_syn_reg_5_ ( .D(ptr_w_syn_1[5]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[5]) );
  DFFR_X1 ptr_w_syn_reg_4_ ( .D(ptr_w_syn_1[4]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[4]) );
  DFFR_X1 ptr_w_syn_reg_3_ ( .D(ptr_w_syn_1[3]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[3]) );
  DFFR_X1 ptr_w_syn_reg_2_ ( .D(ptr_w_syn_1[2]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[2]) );
  DFFR_X1 ptr_w_syn_reg_1_ ( .D(ptr_w_syn_1[1]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[1]), .QN(n32) );
  DFFR_X1 ptr_w_syn_reg_0_ ( .D(ptr_w_syn_1[0]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn[0]) );
  DFFR_X1 ptr_r_syn_reg_8_ ( .D(ptr_r_syn_1[8]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[8]) );
  DFFR_X1 ptr_r_syn_reg_7_ ( .D(ptr_r_syn_1[7]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[7]) );
  DFFR_X1 ptr_r_syn_reg_6_ ( .D(ptr_r_syn_1[6]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[6]) );
  DFFR_X1 ptr_r_syn_reg_5_ ( .D(ptr_r_syn_1[5]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[5]) );
  DFFR_X1 ptr_r_syn_reg_4_ ( .D(ptr_r_syn_1[4]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[4]) );
  DFFR_X1 ptr_r_syn_reg_3_ ( .D(ptr_r_syn_1[3]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[3]) );
  DFFR_X1 ptr_r_syn_reg_2_ ( .D(ptr_r_syn_1[2]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[2]) );
  DFFR_X1 ptr_r_syn_reg_1_ ( .D(ptr_r_syn_1[1]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[1]), .QN(n16) );
  DFFR_X1 ptr_r_syn_reg_0_ ( .D(ptr_r_syn_1[0]), .CK(w_clk), .RN(reset_n), 
        .QN(n17) );
  DFFR_X1 ptr_r_syn_1_reg_8_ ( .D(ptr_r[8]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[8]) );
  DFFR_X1 ptr_w_syn_1_reg_8_ ( .D(ptr_w[8]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[8]) );
  DFFR_X1 ptr_r_syn_1_reg_4_ ( .D(ptr_r[4]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[4]) );
  DFFR_X1 ptr_w_syn_1_reg_7_ ( .D(ptr_w[7]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[7]) );
  DFFR_X1 ptr_r_syn_1_reg_7_ ( .D(ptr_r[7]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[7]) );
  DFFR_X1 ptr_r_syn_1_reg_5_ ( .D(ptr_r[5]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[5]) );
  DFFR_X1 ptr_w_syn_1_reg_5_ ( .D(ptr_w[5]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[5]) );
  DFFR_X1 ptr_w_syn_1_reg_6_ ( .D(ptr_w[6]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[6]) );
  DFFR_X1 ptr_w_syn_1_reg_4_ ( .D(ptr_w[4]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[4]) );
  DFFR_X1 ptr_w_syn_1_reg_3_ ( .D(ptr_w[3]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[3]) );
  DFFR_X1 ptr_w_syn_1_reg_2_ ( .D(ptr_w[2]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[2]) );
  DFFR_X1 ptr_r_syn_1_reg_2_ ( .D(ptr_r[2]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[2]) );
  DFFR_X1 ptr_w_syn_1_reg_0_ ( .D(ptr_w[0]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[0]) );
  DFFR_X1 ptr_r_syn_1_reg_0_ ( .D(ptr_r[0]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[0]) );
  DFFR_X1 ptr_w_syn_1_reg_1_ ( .D(ptr_w[1]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[1]) );
  DFFR_X1 ptr_r_syn_1_reg_1_ ( .D(ptr_r[1]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[1]) );
  DFFR_X1 ptr_r_syn_1_reg_3_ ( .D(ptr_r[3]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[3]) );
  DFFR_X1 ptr_r_syn_1_reg_6_ ( .D(ptr_r[6]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[6]) );
  INV_X1 U3 ( .A(rd), .ZN(n34) );
  INV_X1 U5 ( .A(n3), .ZN(full) );
  AND2_X1 U6 ( .A1(wr), .A2(n3), .ZN(we_enable) );
  NAND3_X1 U7 ( .A1(n40), .A2(n5), .A3(N4), .ZN(n3) );
  INV_X1 U10 ( .A(ptr_w[1]), .ZN(n18) );
  INV_X1 U11 ( .A(ptr_r[0]), .ZN(n1) );
  INV_X1 U12 ( .A(ptr_r[1]), .ZN(n2) );
  XNOR2_X1 U13 ( .A(ptr_r_syn[3]), .B(ptr_w[3]), .ZN(n11) );
  XNOR2_X1 U14 ( .A(ptr_r_syn[2]), .B(ptr_w[2]), .ZN(n10) );
  NOR2_X1 U15 ( .A1(n17), .A2(ptr_w[0]), .ZN(n6) );
  OAI22_X1 U16 ( .A1(n6), .A2(n18), .B1(ptr_r_syn[1]), .B2(n6), .ZN(n9) );
  AND2_X1 U17 ( .A1(ptr_w[0]), .A2(n17), .ZN(n7) );
  OAI22_X1 U18 ( .A1(ptr_w[1]), .A2(n7), .B1(n7), .B2(n16), .ZN(n8) );
  NAND4_X1 U19 ( .A1(n11), .A2(n10), .A3(n9), .A4(n8), .ZN(n15) );
  XOR2_X1 U20 ( .A(ptr_r_syn[6]), .B(ptr_w[6]), .Z(n14) );
  XOR2_X1 U21 ( .A(ptr_r_syn[4]), .B(ptr_w[4]), .Z(n13) );
  XOR2_X1 U22 ( .A(ptr_r_syn[5]), .B(ptr_w[5]), .Z(n12) );
  NOR4_X1 U23 ( .A1(n15), .A2(n14), .A3(n13), .A4(n12), .ZN(N4) );
  XNOR2_X1 U24 ( .A(ptr_r[8]), .B(ptr_w_syn[8]), .ZN(n22) );
  XNOR2_X1 U25 ( .A(ptr_r[7]), .B(ptr_w_syn[7]), .ZN(n21) );
  XNOR2_X1 U26 ( .A(ptr_r[6]), .B(ptr_w_syn[6]), .ZN(n20) );
  XNOR2_X1 U27 ( .A(ptr_r[5]), .B(ptr_w_syn[5]), .ZN(n19) );
  NAND4_X1 U28 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n31) );
  NOR2_X1 U29 ( .A1(n1), .A2(ptr_w_syn[0]), .ZN(n23) );
  OAI22_X1 U30 ( .A1(n23), .A2(n32), .B1(ptr_r[1]), .B2(n23), .ZN(n27) );
  AND2_X1 U31 ( .A1(ptr_w_syn[0]), .A2(n1), .ZN(n24) );
  OAI22_X1 U32 ( .A1(ptr_w_syn[1]), .A2(n24), .B1(n24), .B2(n2), .ZN(n26) );
  XNOR2_X1 U33 ( .A(ptr_r[2]), .B(ptr_w_syn[2]), .ZN(n25) );
  NAND3_X1 U34 ( .A1(n27), .A2(n26), .A3(n25), .ZN(n30) );
  XOR2_X1 U35 ( .A(ptr_r[3]), .B(ptr_w_syn[3]), .Z(n29) );
  XOR2_X1 U36 ( .A(ptr_r[4]), .B(ptr_w_syn[4]), .Z(n28) );
  NOR4_X1 U37 ( .A1(n31), .A2(n30), .A3(n29), .A4(n28), .ZN(empty) );
endmodule


module reg_memory_file_addr_size8_word_width8_1 ( we_s, clk, addr_r, addr_w, 
        data_w, data_r );
  input [7:0] addr_r;
  input [7:0] addr_w;
  input [7:0] data_w;
  output [7:0] data_r;
  input we_s, clk;
  wire   n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095;
  wire   [2047:0] reg_mem;

  DFF_X1 reg_mem_reg_0__7_ ( .D(n7944), .CK(clk), .Q(reg_mem[2047]) );
  DFF_X1 reg_mem_reg_0__6_ ( .D(n7943), .CK(clk), .Q(reg_mem[2046]) );
  DFF_X1 reg_mem_reg_0__5_ ( .D(n7942), .CK(clk), .Q(reg_mem[2045]) );
  DFF_X1 reg_mem_reg_0__4_ ( .D(n7941), .CK(clk), .Q(reg_mem[2044]) );
  DFF_X1 reg_mem_reg_0__3_ ( .D(n7940), .CK(clk), .Q(reg_mem[2043]) );
  DFF_X1 reg_mem_reg_0__2_ ( .D(n7939), .CK(clk), .Q(reg_mem[2042]) );
  DFF_X1 reg_mem_reg_0__1_ ( .D(n7938), .CK(clk), .Q(reg_mem[2041]) );
  DFF_X1 reg_mem_reg_0__0_ ( .D(n7937), .CK(clk), .Q(reg_mem[2040]) );
  DFF_X1 reg_mem_reg_1__7_ ( .D(n7367), .CK(clk), .Q(reg_mem[2039]) );
  DFF_X1 reg_mem_reg_1__6_ ( .D(n7366), .CK(clk), .Q(reg_mem[2038]) );
  DFF_X1 reg_mem_reg_1__5_ ( .D(n7365), .CK(clk), .Q(reg_mem[2037]) );
  DFF_X1 reg_mem_reg_1__4_ ( .D(n7364), .CK(clk), .Q(reg_mem[2036]) );
  DFF_X1 reg_mem_reg_1__3_ ( .D(n7363), .CK(clk), .Q(reg_mem[2035]) );
  DFF_X1 reg_mem_reg_1__2_ ( .D(n7362), .CK(clk), .Q(reg_mem[2034]) );
  DFF_X1 reg_mem_reg_1__1_ ( .D(n7361), .CK(clk), .Q(reg_mem[2033]) );
  DFF_X1 reg_mem_reg_1__0_ ( .D(n7360), .CK(clk), .Q(reg_mem[2032]) );
  DFF_X1 reg_mem_reg_2__7_ ( .D(n8520), .CK(clk), .Q(reg_mem[2031]) );
  DFF_X1 reg_mem_reg_2__6_ ( .D(n8519), .CK(clk), .Q(reg_mem[2030]) );
  DFF_X1 reg_mem_reg_2__5_ ( .D(n8518), .CK(clk), .Q(reg_mem[2029]) );
  DFF_X1 reg_mem_reg_2__4_ ( .D(n8517), .CK(clk), .Q(reg_mem[2028]) );
  DFF_X1 reg_mem_reg_2__3_ ( .D(n8516), .CK(clk), .Q(reg_mem[2027]) );
  DFF_X1 reg_mem_reg_2__2_ ( .D(n8515), .CK(clk), .Q(reg_mem[2026]) );
  DFF_X1 reg_mem_reg_2__1_ ( .D(n8514), .CK(clk), .Q(reg_mem[2025]) );
  DFF_X1 reg_mem_reg_2__0_ ( .D(n8513), .CK(clk), .Q(reg_mem[2024]) );
  DFF_X1 reg_mem_reg_3__7_ ( .D(n6791), .CK(clk), .Q(reg_mem[2023]) );
  DFF_X1 reg_mem_reg_3__6_ ( .D(n6790), .CK(clk), .Q(reg_mem[2022]) );
  DFF_X1 reg_mem_reg_3__5_ ( .D(n6789), .CK(clk), .Q(reg_mem[2021]) );
  DFF_X1 reg_mem_reg_3__4_ ( .D(n6788), .CK(clk), .Q(reg_mem[2020]) );
  DFF_X1 reg_mem_reg_3__3_ ( .D(n6787), .CK(clk), .Q(reg_mem[2019]) );
  DFF_X1 reg_mem_reg_3__2_ ( .D(n6786), .CK(clk), .Q(reg_mem[2018]) );
  DFF_X1 reg_mem_reg_3__1_ ( .D(n6785), .CK(clk), .Q(reg_mem[2017]) );
  DFF_X1 reg_mem_reg_3__0_ ( .D(n6784), .CK(clk), .Q(reg_mem[2016]) );
  DFF_X1 reg_mem_reg_4__7_ ( .D(n8088), .CK(clk), .Q(reg_mem[2015]) );
  DFF_X1 reg_mem_reg_4__6_ ( .D(n8087), .CK(clk), .Q(reg_mem[2014]) );
  DFF_X1 reg_mem_reg_4__5_ ( .D(n8086), .CK(clk), .Q(reg_mem[2013]) );
  DFF_X1 reg_mem_reg_4__4_ ( .D(n8085), .CK(clk), .Q(reg_mem[2012]) );
  DFF_X1 reg_mem_reg_4__3_ ( .D(n8084), .CK(clk), .Q(reg_mem[2011]) );
  DFF_X1 reg_mem_reg_4__2_ ( .D(n8083), .CK(clk), .Q(reg_mem[2010]) );
  DFF_X1 reg_mem_reg_4__1_ ( .D(n8082), .CK(clk), .Q(reg_mem[2009]) );
  DFF_X1 reg_mem_reg_4__0_ ( .D(n8081), .CK(clk), .Q(reg_mem[2008]) );
  DFF_X1 reg_mem_reg_5__7_ ( .D(n7511), .CK(clk), .Q(reg_mem[2007]) );
  DFF_X1 reg_mem_reg_5__6_ ( .D(n7510), .CK(clk), .Q(reg_mem[2006]) );
  DFF_X1 reg_mem_reg_5__5_ ( .D(n7509), .CK(clk), .Q(reg_mem[2005]) );
  DFF_X1 reg_mem_reg_5__4_ ( .D(n7508), .CK(clk), .Q(reg_mem[2004]) );
  DFF_X1 reg_mem_reg_5__3_ ( .D(n7507), .CK(clk), .Q(reg_mem[2003]) );
  DFF_X1 reg_mem_reg_5__2_ ( .D(n7506), .CK(clk), .Q(reg_mem[2002]) );
  DFF_X1 reg_mem_reg_5__1_ ( .D(n7505), .CK(clk), .Q(reg_mem[2001]) );
  DFF_X1 reg_mem_reg_5__0_ ( .D(n7504), .CK(clk), .Q(reg_mem[2000]) );
  DFF_X1 reg_mem_reg_6__7_ ( .D(n8664), .CK(clk), .Q(reg_mem[1999]) );
  DFF_X1 reg_mem_reg_6__6_ ( .D(n8663), .CK(clk), .Q(reg_mem[1998]) );
  DFF_X1 reg_mem_reg_6__5_ ( .D(n8662), .CK(clk), .Q(reg_mem[1997]) );
  DFF_X1 reg_mem_reg_6__4_ ( .D(n8661), .CK(clk), .Q(reg_mem[1996]) );
  DFF_X1 reg_mem_reg_6__3_ ( .D(n8660), .CK(clk), .Q(reg_mem[1995]) );
  DFF_X1 reg_mem_reg_6__2_ ( .D(n8659), .CK(clk), .Q(reg_mem[1994]) );
  DFF_X1 reg_mem_reg_6__1_ ( .D(n8658), .CK(clk), .Q(reg_mem[1993]) );
  DFF_X1 reg_mem_reg_6__0_ ( .D(n8657), .CK(clk), .Q(reg_mem[1992]) );
  DFF_X1 reg_mem_reg_7__7_ ( .D(n6935), .CK(clk), .Q(reg_mem[1991]) );
  DFF_X1 reg_mem_reg_7__6_ ( .D(n6934), .CK(clk), .Q(reg_mem[1990]) );
  DFF_X1 reg_mem_reg_7__5_ ( .D(n6933), .CK(clk), .Q(reg_mem[1989]) );
  DFF_X1 reg_mem_reg_7__4_ ( .D(n6932), .CK(clk), .Q(reg_mem[1988]) );
  DFF_X1 reg_mem_reg_7__3_ ( .D(n6931), .CK(clk), .Q(reg_mem[1987]) );
  DFF_X1 reg_mem_reg_7__2_ ( .D(n6930), .CK(clk), .Q(reg_mem[1986]) );
  DFF_X1 reg_mem_reg_7__1_ ( .D(n6929), .CK(clk), .Q(reg_mem[1985]) );
  DFF_X1 reg_mem_reg_7__0_ ( .D(n6928), .CK(clk), .Q(reg_mem[1984]) );
  DFF_X1 reg_mem_reg_8__7_ ( .D(n8232), .CK(clk), .Q(reg_mem[1983]) );
  DFF_X1 reg_mem_reg_8__6_ ( .D(n8231), .CK(clk), .Q(reg_mem[1982]) );
  DFF_X1 reg_mem_reg_8__5_ ( .D(n8230), .CK(clk), .Q(reg_mem[1981]) );
  DFF_X1 reg_mem_reg_8__4_ ( .D(n8229), .CK(clk), .Q(reg_mem[1980]) );
  DFF_X1 reg_mem_reg_8__3_ ( .D(n8228), .CK(clk), .Q(reg_mem[1979]) );
  DFF_X1 reg_mem_reg_8__2_ ( .D(n8227), .CK(clk), .Q(reg_mem[1978]) );
  DFF_X1 reg_mem_reg_8__1_ ( .D(n8226), .CK(clk), .Q(reg_mem[1977]) );
  DFF_X1 reg_mem_reg_8__0_ ( .D(n8225), .CK(clk), .Q(reg_mem[1976]) );
  DFF_X1 reg_mem_reg_9__7_ ( .D(n7655), .CK(clk), .Q(reg_mem[1975]) );
  DFF_X1 reg_mem_reg_9__6_ ( .D(n7654), .CK(clk), .Q(reg_mem[1974]) );
  DFF_X1 reg_mem_reg_9__5_ ( .D(n7653), .CK(clk), .Q(reg_mem[1973]) );
  DFF_X1 reg_mem_reg_9__4_ ( .D(n7652), .CK(clk), .Q(reg_mem[1972]) );
  DFF_X1 reg_mem_reg_9__3_ ( .D(n7651), .CK(clk), .Q(reg_mem[1971]) );
  DFF_X1 reg_mem_reg_9__2_ ( .D(n7650), .CK(clk), .Q(reg_mem[1970]) );
  DFF_X1 reg_mem_reg_9__1_ ( .D(n7649), .CK(clk), .Q(reg_mem[1969]) );
  DFF_X1 reg_mem_reg_9__0_ ( .D(n7648), .CK(clk), .Q(reg_mem[1968]) );
  DFF_X1 reg_mem_reg_10__7_ ( .D(n8808), .CK(clk), .Q(reg_mem[1967]) );
  DFF_X1 reg_mem_reg_10__6_ ( .D(n8807), .CK(clk), .Q(reg_mem[1966]) );
  DFF_X1 reg_mem_reg_10__5_ ( .D(n8806), .CK(clk), .Q(reg_mem[1965]) );
  DFF_X1 reg_mem_reg_10__4_ ( .D(n8805), .CK(clk), .Q(reg_mem[1964]) );
  DFF_X1 reg_mem_reg_10__3_ ( .D(n8804), .CK(clk), .Q(reg_mem[1963]) );
  DFF_X1 reg_mem_reg_10__2_ ( .D(n8803), .CK(clk), .Q(reg_mem[1962]) );
  DFF_X1 reg_mem_reg_10__1_ ( .D(n8802), .CK(clk), .Q(reg_mem[1961]) );
  DFF_X1 reg_mem_reg_10__0_ ( .D(n8801), .CK(clk), .Q(reg_mem[1960]) );
  DFF_X1 reg_mem_reg_11__7_ ( .D(n7079), .CK(clk), .Q(reg_mem[1959]) );
  DFF_X1 reg_mem_reg_11__6_ ( .D(n7078), .CK(clk), .Q(reg_mem[1958]) );
  DFF_X1 reg_mem_reg_11__5_ ( .D(n7077), .CK(clk), .Q(reg_mem[1957]) );
  DFF_X1 reg_mem_reg_11__4_ ( .D(n7076), .CK(clk), .Q(reg_mem[1956]) );
  DFF_X1 reg_mem_reg_11__3_ ( .D(n7075), .CK(clk), .Q(reg_mem[1955]) );
  DFF_X1 reg_mem_reg_11__2_ ( .D(n7074), .CK(clk), .Q(reg_mem[1954]) );
  DFF_X1 reg_mem_reg_11__1_ ( .D(n7073), .CK(clk), .Q(reg_mem[1953]) );
  DFF_X1 reg_mem_reg_11__0_ ( .D(n7072), .CK(clk), .Q(reg_mem[1952]) );
  DFF_X1 reg_mem_reg_12__7_ ( .D(n8376), .CK(clk), .Q(reg_mem[1951]) );
  DFF_X1 reg_mem_reg_12__6_ ( .D(n8375), .CK(clk), .Q(reg_mem[1950]) );
  DFF_X1 reg_mem_reg_12__5_ ( .D(n8374), .CK(clk), .Q(reg_mem[1949]) );
  DFF_X1 reg_mem_reg_12__4_ ( .D(n8373), .CK(clk), .Q(reg_mem[1948]) );
  DFF_X1 reg_mem_reg_12__3_ ( .D(n8372), .CK(clk), .Q(reg_mem[1947]) );
  DFF_X1 reg_mem_reg_12__2_ ( .D(n8371), .CK(clk), .Q(reg_mem[1946]) );
  DFF_X1 reg_mem_reg_12__1_ ( .D(n8370), .CK(clk), .Q(reg_mem[1945]) );
  DFF_X1 reg_mem_reg_12__0_ ( .D(n8369), .CK(clk), .Q(reg_mem[1944]) );
  DFF_X1 reg_mem_reg_13__7_ ( .D(n7799), .CK(clk), .Q(reg_mem[1943]) );
  DFF_X1 reg_mem_reg_13__6_ ( .D(n7798), .CK(clk), .Q(reg_mem[1942]) );
  DFF_X1 reg_mem_reg_13__5_ ( .D(n7797), .CK(clk), .Q(reg_mem[1941]) );
  DFF_X1 reg_mem_reg_13__4_ ( .D(n7796), .CK(clk), .Q(reg_mem[1940]) );
  DFF_X1 reg_mem_reg_13__3_ ( .D(n7795), .CK(clk), .Q(reg_mem[1939]) );
  DFF_X1 reg_mem_reg_13__2_ ( .D(n7794), .CK(clk), .Q(reg_mem[1938]) );
  DFF_X1 reg_mem_reg_13__1_ ( .D(n7793), .CK(clk), .Q(reg_mem[1937]) );
  DFF_X1 reg_mem_reg_13__0_ ( .D(n7792), .CK(clk), .Q(reg_mem[1936]) );
  DFF_X1 reg_mem_reg_14__7_ ( .D(n8952), .CK(clk), .Q(reg_mem[1935]) );
  DFF_X1 reg_mem_reg_14__6_ ( .D(n8951), .CK(clk), .Q(reg_mem[1934]) );
  DFF_X1 reg_mem_reg_14__5_ ( .D(n8950), .CK(clk), .Q(reg_mem[1933]) );
  DFF_X1 reg_mem_reg_14__4_ ( .D(n8949), .CK(clk), .Q(reg_mem[1932]) );
  DFF_X1 reg_mem_reg_14__3_ ( .D(n8948), .CK(clk), .Q(reg_mem[1931]) );
  DFF_X1 reg_mem_reg_14__2_ ( .D(n8947), .CK(clk), .Q(reg_mem[1930]) );
  DFF_X1 reg_mem_reg_14__1_ ( .D(n8946), .CK(clk), .Q(reg_mem[1929]) );
  DFF_X1 reg_mem_reg_14__0_ ( .D(n8945), .CK(clk), .Q(reg_mem[1928]) );
  DFF_X1 reg_mem_reg_15__7_ ( .D(n7223), .CK(clk), .Q(reg_mem[1927]) );
  DFF_X1 reg_mem_reg_15__6_ ( .D(n7222), .CK(clk), .Q(reg_mem[1926]) );
  DFF_X1 reg_mem_reg_15__5_ ( .D(n7221), .CK(clk), .Q(reg_mem[1925]) );
  DFF_X1 reg_mem_reg_15__4_ ( .D(n7220), .CK(clk), .Q(reg_mem[1924]) );
  DFF_X1 reg_mem_reg_15__3_ ( .D(n7219), .CK(clk), .Q(reg_mem[1923]) );
  DFF_X1 reg_mem_reg_15__2_ ( .D(n7218), .CK(clk), .Q(reg_mem[1922]) );
  DFF_X1 reg_mem_reg_15__1_ ( .D(n7217), .CK(clk), .Q(reg_mem[1921]) );
  DFF_X1 reg_mem_reg_15__0_ ( .D(n7216), .CK(clk), .Q(reg_mem[1920]) );
  DFF_X1 reg_mem_reg_16__7_ ( .D(n7953), .CK(clk), .Q(reg_mem[1919]) );
  DFF_X1 reg_mem_reg_16__6_ ( .D(n7952), .CK(clk), .Q(reg_mem[1918]) );
  DFF_X1 reg_mem_reg_16__5_ ( .D(n7951), .CK(clk), .Q(reg_mem[1917]) );
  DFF_X1 reg_mem_reg_16__4_ ( .D(n7950), .CK(clk), .Q(reg_mem[1916]) );
  DFF_X1 reg_mem_reg_16__3_ ( .D(n7949), .CK(clk), .Q(reg_mem[1915]) );
  DFF_X1 reg_mem_reg_16__2_ ( .D(n7948), .CK(clk), .Q(reg_mem[1914]) );
  DFF_X1 reg_mem_reg_16__1_ ( .D(n7947), .CK(clk), .Q(reg_mem[1913]) );
  DFF_X1 reg_mem_reg_16__0_ ( .D(n7946), .CK(clk), .Q(reg_mem[1912]) );
  DFF_X1 reg_mem_reg_17__7_ ( .D(n7376), .CK(clk), .Q(reg_mem[1911]) );
  DFF_X1 reg_mem_reg_17__6_ ( .D(n7375), .CK(clk), .Q(reg_mem[1910]) );
  DFF_X1 reg_mem_reg_17__5_ ( .D(n7374), .CK(clk), .Q(reg_mem[1909]) );
  DFF_X1 reg_mem_reg_17__4_ ( .D(n7373), .CK(clk), .Q(reg_mem[1908]) );
  DFF_X1 reg_mem_reg_17__3_ ( .D(n7372), .CK(clk), .Q(reg_mem[1907]) );
  DFF_X1 reg_mem_reg_17__2_ ( .D(n7371), .CK(clk), .Q(reg_mem[1906]) );
  DFF_X1 reg_mem_reg_17__1_ ( .D(n7370), .CK(clk), .Q(reg_mem[1905]) );
  DFF_X1 reg_mem_reg_17__0_ ( .D(n7369), .CK(clk), .Q(reg_mem[1904]) );
  DFF_X1 reg_mem_reg_18__7_ ( .D(n8529), .CK(clk), .Q(reg_mem[1903]) );
  DFF_X1 reg_mem_reg_18__6_ ( .D(n8528), .CK(clk), .Q(reg_mem[1902]) );
  DFF_X1 reg_mem_reg_18__5_ ( .D(n8527), .CK(clk), .Q(reg_mem[1901]) );
  DFF_X1 reg_mem_reg_18__4_ ( .D(n8526), .CK(clk), .Q(reg_mem[1900]) );
  DFF_X1 reg_mem_reg_18__3_ ( .D(n8525), .CK(clk), .Q(reg_mem[1899]) );
  DFF_X1 reg_mem_reg_18__2_ ( .D(n8524), .CK(clk), .Q(reg_mem[1898]) );
  DFF_X1 reg_mem_reg_18__1_ ( .D(n8523), .CK(clk), .Q(reg_mem[1897]) );
  DFF_X1 reg_mem_reg_18__0_ ( .D(n8522), .CK(clk), .Q(reg_mem[1896]) );
  DFF_X1 reg_mem_reg_19__7_ ( .D(n6800), .CK(clk), .Q(reg_mem[1895]) );
  DFF_X1 reg_mem_reg_19__6_ ( .D(n6799), .CK(clk), .Q(reg_mem[1894]) );
  DFF_X1 reg_mem_reg_19__5_ ( .D(n6798), .CK(clk), .Q(reg_mem[1893]) );
  DFF_X1 reg_mem_reg_19__4_ ( .D(n6797), .CK(clk), .Q(reg_mem[1892]) );
  DFF_X1 reg_mem_reg_19__3_ ( .D(n6796), .CK(clk), .Q(reg_mem[1891]) );
  DFF_X1 reg_mem_reg_19__2_ ( .D(n6795), .CK(clk), .Q(reg_mem[1890]) );
  DFF_X1 reg_mem_reg_19__1_ ( .D(n6794), .CK(clk), .Q(reg_mem[1889]) );
  DFF_X1 reg_mem_reg_19__0_ ( .D(n6793), .CK(clk), .Q(reg_mem[1888]) );
  DFF_X1 reg_mem_reg_20__7_ ( .D(n8097), .CK(clk), .Q(reg_mem[1887]) );
  DFF_X1 reg_mem_reg_20__6_ ( .D(n8096), .CK(clk), .Q(reg_mem[1886]) );
  DFF_X1 reg_mem_reg_20__5_ ( .D(n8095), .CK(clk), .Q(reg_mem[1885]) );
  DFF_X1 reg_mem_reg_20__4_ ( .D(n8094), .CK(clk), .Q(reg_mem[1884]) );
  DFF_X1 reg_mem_reg_20__3_ ( .D(n8093), .CK(clk), .Q(reg_mem[1883]) );
  DFF_X1 reg_mem_reg_20__2_ ( .D(n8092), .CK(clk), .Q(reg_mem[1882]) );
  DFF_X1 reg_mem_reg_20__1_ ( .D(n8091), .CK(clk), .Q(reg_mem[1881]) );
  DFF_X1 reg_mem_reg_20__0_ ( .D(n8090), .CK(clk), .Q(reg_mem[1880]) );
  DFF_X1 reg_mem_reg_21__7_ ( .D(n7520), .CK(clk), .Q(reg_mem[1879]) );
  DFF_X1 reg_mem_reg_21__6_ ( .D(n7519), .CK(clk), .Q(reg_mem[1878]) );
  DFF_X1 reg_mem_reg_21__5_ ( .D(n7518), .CK(clk), .Q(reg_mem[1877]) );
  DFF_X1 reg_mem_reg_21__4_ ( .D(n7517), .CK(clk), .Q(reg_mem[1876]) );
  DFF_X1 reg_mem_reg_21__3_ ( .D(n7516), .CK(clk), .Q(reg_mem[1875]) );
  DFF_X1 reg_mem_reg_21__2_ ( .D(n7515), .CK(clk), .Q(reg_mem[1874]) );
  DFF_X1 reg_mem_reg_21__1_ ( .D(n7514), .CK(clk), .Q(reg_mem[1873]) );
  DFF_X1 reg_mem_reg_21__0_ ( .D(n7513), .CK(clk), .Q(reg_mem[1872]) );
  DFF_X1 reg_mem_reg_22__7_ ( .D(n8673), .CK(clk), .Q(reg_mem[1871]) );
  DFF_X1 reg_mem_reg_22__6_ ( .D(n8672), .CK(clk), .Q(reg_mem[1870]) );
  DFF_X1 reg_mem_reg_22__5_ ( .D(n8671), .CK(clk), .Q(reg_mem[1869]) );
  DFF_X1 reg_mem_reg_22__4_ ( .D(n8670), .CK(clk), .Q(reg_mem[1868]) );
  DFF_X1 reg_mem_reg_22__3_ ( .D(n8669), .CK(clk), .Q(reg_mem[1867]) );
  DFF_X1 reg_mem_reg_22__2_ ( .D(n8668), .CK(clk), .Q(reg_mem[1866]) );
  DFF_X1 reg_mem_reg_22__1_ ( .D(n8667), .CK(clk), .Q(reg_mem[1865]) );
  DFF_X1 reg_mem_reg_22__0_ ( .D(n8666), .CK(clk), .Q(reg_mem[1864]) );
  DFF_X1 reg_mem_reg_23__7_ ( .D(n6944), .CK(clk), .Q(reg_mem[1863]) );
  DFF_X1 reg_mem_reg_23__6_ ( .D(n6943), .CK(clk), .Q(reg_mem[1862]) );
  DFF_X1 reg_mem_reg_23__5_ ( .D(n6942), .CK(clk), .Q(reg_mem[1861]) );
  DFF_X1 reg_mem_reg_23__4_ ( .D(n6941), .CK(clk), .Q(reg_mem[1860]) );
  DFF_X1 reg_mem_reg_23__3_ ( .D(n6940), .CK(clk), .Q(reg_mem[1859]) );
  DFF_X1 reg_mem_reg_23__2_ ( .D(n6939), .CK(clk), .Q(reg_mem[1858]) );
  DFF_X1 reg_mem_reg_23__1_ ( .D(n6938), .CK(clk), .Q(reg_mem[1857]) );
  DFF_X1 reg_mem_reg_23__0_ ( .D(n6937), .CK(clk), .Q(reg_mem[1856]) );
  DFF_X1 reg_mem_reg_24__7_ ( .D(n8241), .CK(clk), .Q(reg_mem[1855]) );
  DFF_X1 reg_mem_reg_24__6_ ( .D(n8240), .CK(clk), .Q(reg_mem[1854]) );
  DFF_X1 reg_mem_reg_24__5_ ( .D(n8239), .CK(clk), .Q(reg_mem[1853]) );
  DFF_X1 reg_mem_reg_24__4_ ( .D(n8238), .CK(clk), .Q(reg_mem[1852]) );
  DFF_X1 reg_mem_reg_24__3_ ( .D(n8237), .CK(clk), .Q(reg_mem[1851]) );
  DFF_X1 reg_mem_reg_24__2_ ( .D(n8236), .CK(clk), .Q(reg_mem[1850]) );
  DFF_X1 reg_mem_reg_24__1_ ( .D(n8235), .CK(clk), .Q(reg_mem[1849]) );
  DFF_X1 reg_mem_reg_24__0_ ( .D(n8234), .CK(clk), .Q(reg_mem[1848]) );
  DFF_X1 reg_mem_reg_25__7_ ( .D(n7664), .CK(clk), .Q(reg_mem[1847]) );
  DFF_X1 reg_mem_reg_25__6_ ( .D(n7663), .CK(clk), .Q(reg_mem[1846]) );
  DFF_X1 reg_mem_reg_25__5_ ( .D(n7662), .CK(clk), .Q(reg_mem[1845]) );
  DFF_X1 reg_mem_reg_25__4_ ( .D(n7661), .CK(clk), .Q(reg_mem[1844]) );
  DFF_X1 reg_mem_reg_25__3_ ( .D(n7660), .CK(clk), .Q(reg_mem[1843]) );
  DFF_X1 reg_mem_reg_25__2_ ( .D(n7659), .CK(clk), .Q(reg_mem[1842]) );
  DFF_X1 reg_mem_reg_25__1_ ( .D(n7658), .CK(clk), .Q(reg_mem[1841]) );
  DFF_X1 reg_mem_reg_25__0_ ( .D(n7657), .CK(clk), .Q(reg_mem[1840]) );
  DFF_X1 reg_mem_reg_26__7_ ( .D(n8817), .CK(clk), .Q(reg_mem[1839]) );
  DFF_X1 reg_mem_reg_26__6_ ( .D(n8816), .CK(clk), .Q(reg_mem[1838]) );
  DFF_X1 reg_mem_reg_26__5_ ( .D(n8815), .CK(clk), .Q(reg_mem[1837]) );
  DFF_X1 reg_mem_reg_26__4_ ( .D(n8814), .CK(clk), .Q(reg_mem[1836]) );
  DFF_X1 reg_mem_reg_26__3_ ( .D(n8813), .CK(clk), .Q(reg_mem[1835]) );
  DFF_X1 reg_mem_reg_26__2_ ( .D(n8812), .CK(clk), .Q(reg_mem[1834]) );
  DFF_X1 reg_mem_reg_26__1_ ( .D(n8811), .CK(clk), .Q(reg_mem[1833]) );
  DFF_X1 reg_mem_reg_26__0_ ( .D(n8810), .CK(clk), .Q(reg_mem[1832]) );
  DFF_X1 reg_mem_reg_27__7_ ( .D(n7088), .CK(clk), .Q(reg_mem[1831]) );
  DFF_X1 reg_mem_reg_27__6_ ( .D(n7087), .CK(clk), .Q(reg_mem[1830]) );
  DFF_X1 reg_mem_reg_27__5_ ( .D(n7086), .CK(clk), .Q(reg_mem[1829]) );
  DFF_X1 reg_mem_reg_27__4_ ( .D(n7085), .CK(clk), .Q(reg_mem[1828]) );
  DFF_X1 reg_mem_reg_27__3_ ( .D(n7084), .CK(clk), .Q(reg_mem[1827]) );
  DFF_X1 reg_mem_reg_27__2_ ( .D(n7083), .CK(clk), .Q(reg_mem[1826]) );
  DFF_X1 reg_mem_reg_27__1_ ( .D(n7082), .CK(clk), .Q(reg_mem[1825]) );
  DFF_X1 reg_mem_reg_27__0_ ( .D(n7081), .CK(clk), .Q(reg_mem[1824]) );
  DFF_X1 reg_mem_reg_28__7_ ( .D(n8385), .CK(clk), .Q(reg_mem[1823]) );
  DFF_X1 reg_mem_reg_28__6_ ( .D(n8384), .CK(clk), .Q(reg_mem[1822]) );
  DFF_X1 reg_mem_reg_28__5_ ( .D(n8383), .CK(clk), .Q(reg_mem[1821]) );
  DFF_X1 reg_mem_reg_28__4_ ( .D(n8382), .CK(clk), .Q(reg_mem[1820]) );
  DFF_X1 reg_mem_reg_28__3_ ( .D(n8381), .CK(clk), .Q(reg_mem[1819]) );
  DFF_X1 reg_mem_reg_28__2_ ( .D(n8380), .CK(clk), .Q(reg_mem[1818]) );
  DFF_X1 reg_mem_reg_28__1_ ( .D(n8379), .CK(clk), .Q(reg_mem[1817]) );
  DFF_X1 reg_mem_reg_28__0_ ( .D(n8378), .CK(clk), .Q(reg_mem[1816]) );
  DFF_X1 reg_mem_reg_29__7_ ( .D(n7808), .CK(clk), .Q(reg_mem[1815]) );
  DFF_X1 reg_mem_reg_29__6_ ( .D(n7807), .CK(clk), .Q(reg_mem[1814]) );
  DFF_X1 reg_mem_reg_29__5_ ( .D(n7806), .CK(clk), .Q(reg_mem[1813]) );
  DFF_X1 reg_mem_reg_29__4_ ( .D(n7805), .CK(clk), .Q(reg_mem[1812]) );
  DFF_X1 reg_mem_reg_29__3_ ( .D(n7804), .CK(clk), .Q(reg_mem[1811]) );
  DFF_X1 reg_mem_reg_29__2_ ( .D(n7803), .CK(clk), .Q(reg_mem[1810]) );
  DFF_X1 reg_mem_reg_29__1_ ( .D(n7802), .CK(clk), .Q(reg_mem[1809]) );
  DFF_X1 reg_mem_reg_29__0_ ( .D(n7801), .CK(clk), .Q(reg_mem[1808]) );
  DFF_X1 reg_mem_reg_30__7_ ( .D(n8961), .CK(clk), .Q(reg_mem[1807]) );
  DFF_X1 reg_mem_reg_30__6_ ( .D(n8960), .CK(clk), .Q(reg_mem[1806]) );
  DFF_X1 reg_mem_reg_30__5_ ( .D(n8959), .CK(clk), .Q(reg_mem[1805]) );
  DFF_X1 reg_mem_reg_30__4_ ( .D(n8958), .CK(clk), .Q(reg_mem[1804]) );
  DFF_X1 reg_mem_reg_30__3_ ( .D(n8957), .CK(clk), .Q(reg_mem[1803]) );
  DFF_X1 reg_mem_reg_30__2_ ( .D(n8956), .CK(clk), .Q(reg_mem[1802]) );
  DFF_X1 reg_mem_reg_30__1_ ( .D(n8955), .CK(clk), .Q(reg_mem[1801]) );
  DFF_X1 reg_mem_reg_30__0_ ( .D(n8954), .CK(clk), .Q(reg_mem[1800]) );
  DFF_X1 reg_mem_reg_31__7_ ( .D(n7232), .CK(clk), .Q(reg_mem[1799]) );
  DFF_X1 reg_mem_reg_31__6_ ( .D(n7231), .CK(clk), .Q(reg_mem[1798]) );
  DFF_X1 reg_mem_reg_31__5_ ( .D(n7230), .CK(clk), .Q(reg_mem[1797]) );
  DFF_X1 reg_mem_reg_31__4_ ( .D(n7229), .CK(clk), .Q(reg_mem[1796]) );
  DFF_X1 reg_mem_reg_31__3_ ( .D(n7228), .CK(clk), .Q(reg_mem[1795]) );
  DFF_X1 reg_mem_reg_31__2_ ( .D(n7227), .CK(clk), .Q(reg_mem[1794]) );
  DFF_X1 reg_mem_reg_31__1_ ( .D(n7226), .CK(clk), .Q(reg_mem[1793]) );
  DFF_X1 reg_mem_reg_31__0_ ( .D(n7225), .CK(clk), .Q(reg_mem[1792]) );
  DFF_X1 reg_mem_reg_32__7_ ( .D(n7962), .CK(clk), .Q(reg_mem[1791]) );
  DFF_X1 reg_mem_reg_32__6_ ( .D(n7961), .CK(clk), .Q(reg_mem[1790]) );
  DFF_X1 reg_mem_reg_32__5_ ( .D(n7960), .CK(clk), .Q(reg_mem[1789]) );
  DFF_X1 reg_mem_reg_32__4_ ( .D(n7959), .CK(clk), .Q(reg_mem[1788]) );
  DFF_X1 reg_mem_reg_32__3_ ( .D(n7958), .CK(clk), .Q(reg_mem[1787]) );
  DFF_X1 reg_mem_reg_32__2_ ( .D(n7957), .CK(clk), .Q(reg_mem[1786]) );
  DFF_X1 reg_mem_reg_32__1_ ( .D(n7956), .CK(clk), .Q(reg_mem[1785]) );
  DFF_X1 reg_mem_reg_32__0_ ( .D(n7955), .CK(clk), .Q(reg_mem[1784]) );
  DFF_X1 reg_mem_reg_33__7_ ( .D(n7385), .CK(clk), .Q(reg_mem[1783]) );
  DFF_X1 reg_mem_reg_33__6_ ( .D(n7384), .CK(clk), .Q(reg_mem[1782]) );
  DFF_X1 reg_mem_reg_33__5_ ( .D(n7383), .CK(clk), .Q(reg_mem[1781]) );
  DFF_X1 reg_mem_reg_33__4_ ( .D(n7382), .CK(clk), .Q(reg_mem[1780]) );
  DFF_X1 reg_mem_reg_33__3_ ( .D(n7381), .CK(clk), .Q(reg_mem[1779]) );
  DFF_X1 reg_mem_reg_33__2_ ( .D(n7380), .CK(clk), .Q(reg_mem[1778]) );
  DFF_X1 reg_mem_reg_33__1_ ( .D(n7379), .CK(clk), .Q(reg_mem[1777]) );
  DFF_X1 reg_mem_reg_33__0_ ( .D(n7378), .CK(clk), .Q(reg_mem[1776]) );
  DFF_X1 reg_mem_reg_34__7_ ( .D(n8538), .CK(clk), .Q(reg_mem[1775]) );
  DFF_X1 reg_mem_reg_34__6_ ( .D(n8537), .CK(clk), .Q(reg_mem[1774]) );
  DFF_X1 reg_mem_reg_34__5_ ( .D(n8536), .CK(clk), .Q(reg_mem[1773]) );
  DFF_X1 reg_mem_reg_34__4_ ( .D(n8535), .CK(clk), .Q(reg_mem[1772]) );
  DFF_X1 reg_mem_reg_34__3_ ( .D(n8534), .CK(clk), .Q(reg_mem[1771]) );
  DFF_X1 reg_mem_reg_34__2_ ( .D(n8533), .CK(clk), .Q(reg_mem[1770]) );
  DFF_X1 reg_mem_reg_34__1_ ( .D(n8532), .CK(clk), .Q(reg_mem[1769]) );
  DFF_X1 reg_mem_reg_34__0_ ( .D(n8531), .CK(clk), .Q(reg_mem[1768]) );
  DFF_X1 reg_mem_reg_35__7_ ( .D(n6809), .CK(clk), .Q(reg_mem[1767]) );
  DFF_X1 reg_mem_reg_35__6_ ( .D(n6808), .CK(clk), .Q(reg_mem[1766]) );
  DFF_X1 reg_mem_reg_35__5_ ( .D(n6807), .CK(clk), .Q(reg_mem[1765]) );
  DFF_X1 reg_mem_reg_35__4_ ( .D(n6806), .CK(clk), .Q(reg_mem[1764]) );
  DFF_X1 reg_mem_reg_35__3_ ( .D(n6805), .CK(clk), .Q(reg_mem[1763]) );
  DFF_X1 reg_mem_reg_35__2_ ( .D(n6804), .CK(clk), .Q(reg_mem[1762]) );
  DFF_X1 reg_mem_reg_35__1_ ( .D(n6803), .CK(clk), .Q(reg_mem[1761]) );
  DFF_X1 reg_mem_reg_35__0_ ( .D(n6802), .CK(clk), .Q(reg_mem[1760]) );
  DFF_X1 reg_mem_reg_36__7_ ( .D(n8106), .CK(clk), .Q(reg_mem[1759]) );
  DFF_X1 reg_mem_reg_36__6_ ( .D(n8105), .CK(clk), .Q(reg_mem[1758]) );
  DFF_X1 reg_mem_reg_36__5_ ( .D(n8104), .CK(clk), .Q(reg_mem[1757]) );
  DFF_X1 reg_mem_reg_36__4_ ( .D(n8103), .CK(clk), .Q(reg_mem[1756]) );
  DFF_X1 reg_mem_reg_36__3_ ( .D(n8102), .CK(clk), .Q(reg_mem[1755]) );
  DFF_X1 reg_mem_reg_36__2_ ( .D(n8101), .CK(clk), .Q(reg_mem[1754]) );
  DFF_X1 reg_mem_reg_36__1_ ( .D(n8100), .CK(clk), .Q(reg_mem[1753]) );
  DFF_X1 reg_mem_reg_36__0_ ( .D(n8099), .CK(clk), .Q(reg_mem[1752]) );
  DFF_X1 reg_mem_reg_37__7_ ( .D(n7529), .CK(clk), .Q(reg_mem[1751]) );
  DFF_X1 reg_mem_reg_37__6_ ( .D(n7528), .CK(clk), .Q(reg_mem[1750]) );
  DFF_X1 reg_mem_reg_37__5_ ( .D(n7527), .CK(clk), .Q(reg_mem[1749]) );
  DFF_X1 reg_mem_reg_37__4_ ( .D(n7526), .CK(clk), .Q(reg_mem[1748]) );
  DFF_X1 reg_mem_reg_37__3_ ( .D(n7525), .CK(clk), .Q(reg_mem[1747]) );
  DFF_X1 reg_mem_reg_37__2_ ( .D(n7524), .CK(clk), .Q(reg_mem[1746]) );
  DFF_X1 reg_mem_reg_37__1_ ( .D(n7523), .CK(clk), .Q(reg_mem[1745]) );
  DFF_X1 reg_mem_reg_37__0_ ( .D(n7522), .CK(clk), .Q(reg_mem[1744]) );
  DFF_X1 reg_mem_reg_38__7_ ( .D(n8682), .CK(clk), .Q(reg_mem[1743]) );
  DFF_X1 reg_mem_reg_38__6_ ( .D(n8681), .CK(clk), .Q(reg_mem[1742]) );
  DFF_X1 reg_mem_reg_38__5_ ( .D(n8680), .CK(clk), .Q(reg_mem[1741]) );
  DFF_X1 reg_mem_reg_38__4_ ( .D(n8679), .CK(clk), .Q(reg_mem[1740]) );
  DFF_X1 reg_mem_reg_38__3_ ( .D(n8678), .CK(clk), .Q(reg_mem[1739]) );
  DFF_X1 reg_mem_reg_38__2_ ( .D(n8677), .CK(clk), .Q(reg_mem[1738]) );
  DFF_X1 reg_mem_reg_38__1_ ( .D(n8676), .CK(clk), .Q(reg_mem[1737]) );
  DFF_X1 reg_mem_reg_38__0_ ( .D(n8675), .CK(clk), .Q(reg_mem[1736]) );
  DFF_X1 reg_mem_reg_39__7_ ( .D(n6953), .CK(clk), .Q(reg_mem[1735]) );
  DFF_X1 reg_mem_reg_39__6_ ( .D(n6952), .CK(clk), .Q(reg_mem[1734]) );
  DFF_X1 reg_mem_reg_39__5_ ( .D(n6951), .CK(clk), .Q(reg_mem[1733]) );
  DFF_X1 reg_mem_reg_39__4_ ( .D(n6950), .CK(clk), .Q(reg_mem[1732]) );
  DFF_X1 reg_mem_reg_39__3_ ( .D(n6949), .CK(clk), .Q(reg_mem[1731]) );
  DFF_X1 reg_mem_reg_39__2_ ( .D(n6948), .CK(clk), .Q(reg_mem[1730]) );
  DFF_X1 reg_mem_reg_39__1_ ( .D(n6947), .CK(clk), .Q(reg_mem[1729]) );
  DFF_X1 reg_mem_reg_39__0_ ( .D(n6946), .CK(clk), .Q(reg_mem[1728]) );
  DFF_X1 reg_mem_reg_40__7_ ( .D(n8250), .CK(clk), .Q(reg_mem[1727]) );
  DFF_X1 reg_mem_reg_40__6_ ( .D(n8249), .CK(clk), .Q(reg_mem[1726]) );
  DFF_X1 reg_mem_reg_40__5_ ( .D(n8248), .CK(clk), .Q(reg_mem[1725]) );
  DFF_X1 reg_mem_reg_40__4_ ( .D(n8247), .CK(clk), .Q(reg_mem[1724]) );
  DFF_X1 reg_mem_reg_40__3_ ( .D(n8246), .CK(clk), .Q(reg_mem[1723]) );
  DFF_X1 reg_mem_reg_40__2_ ( .D(n8245), .CK(clk), .Q(reg_mem[1722]) );
  DFF_X1 reg_mem_reg_40__1_ ( .D(n8244), .CK(clk), .Q(reg_mem[1721]) );
  DFF_X1 reg_mem_reg_40__0_ ( .D(n8243), .CK(clk), .Q(reg_mem[1720]) );
  DFF_X1 reg_mem_reg_41__7_ ( .D(n7673), .CK(clk), .Q(reg_mem[1719]) );
  DFF_X1 reg_mem_reg_41__6_ ( .D(n7672), .CK(clk), .Q(reg_mem[1718]) );
  DFF_X1 reg_mem_reg_41__5_ ( .D(n7671), .CK(clk), .Q(reg_mem[1717]) );
  DFF_X1 reg_mem_reg_41__4_ ( .D(n7670), .CK(clk), .Q(reg_mem[1716]) );
  DFF_X1 reg_mem_reg_41__3_ ( .D(n7669), .CK(clk), .Q(reg_mem[1715]) );
  DFF_X1 reg_mem_reg_41__2_ ( .D(n7668), .CK(clk), .Q(reg_mem[1714]) );
  DFF_X1 reg_mem_reg_41__1_ ( .D(n7667), .CK(clk), .Q(reg_mem[1713]) );
  DFF_X1 reg_mem_reg_41__0_ ( .D(n7666), .CK(clk), .Q(reg_mem[1712]) );
  DFF_X1 reg_mem_reg_42__7_ ( .D(n8826), .CK(clk), .Q(reg_mem[1711]) );
  DFF_X1 reg_mem_reg_42__6_ ( .D(n8825), .CK(clk), .Q(reg_mem[1710]) );
  DFF_X1 reg_mem_reg_42__5_ ( .D(n8824), .CK(clk), .Q(reg_mem[1709]) );
  DFF_X1 reg_mem_reg_42__4_ ( .D(n8823), .CK(clk), .Q(reg_mem[1708]) );
  DFF_X1 reg_mem_reg_42__3_ ( .D(n8822), .CK(clk), .Q(reg_mem[1707]) );
  DFF_X1 reg_mem_reg_42__2_ ( .D(n8821), .CK(clk), .Q(reg_mem[1706]) );
  DFF_X1 reg_mem_reg_42__1_ ( .D(n8820), .CK(clk), .Q(reg_mem[1705]) );
  DFF_X1 reg_mem_reg_42__0_ ( .D(n8819), .CK(clk), .Q(reg_mem[1704]) );
  DFF_X1 reg_mem_reg_43__7_ ( .D(n7097), .CK(clk), .Q(reg_mem[1703]) );
  DFF_X1 reg_mem_reg_43__6_ ( .D(n7096), .CK(clk), .Q(reg_mem[1702]) );
  DFF_X1 reg_mem_reg_43__5_ ( .D(n7095), .CK(clk), .Q(reg_mem[1701]) );
  DFF_X1 reg_mem_reg_43__4_ ( .D(n7094), .CK(clk), .Q(reg_mem[1700]) );
  DFF_X1 reg_mem_reg_43__3_ ( .D(n7093), .CK(clk), .Q(reg_mem[1699]) );
  DFF_X1 reg_mem_reg_43__2_ ( .D(n7092), .CK(clk), .Q(reg_mem[1698]) );
  DFF_X1 reg_mem_reg_43__1_ ( .D(n7091), .CK(clk), .Q(reg_mem[1697]) );
  DFF_X1 reg_mem_reg_43__0_ ( .D(n7090), .CK(clk), .Q(reg_mem[1696]) );
  DFF_X1 reg_mem_reg_44__7_ ( .D(n8394), .CK(clk), .Q(reg_mem[1695]) );
  DFF_X1 reg_mem_reg_44__6_ ( .D(n8393), .CK(clk), .Q(reg_mem[1694]) );
  DFF_X1 reg_mem_reg_44__5_ ( .D(n8392), .CK(clk), .Q(reg_mem[1693]) );
  DFF_X1 reg_mem_reg_44__4_ ( .D(n8391), .CK(clk), .Q(reg_mem[1692]) );
  DFF_X1 reg_mem_reg_44__3_ ( .D(n8390), .CK(clk), .Q(reg_mem[1691]) );
  DFF_X1 reg_mem_reg_44__2_ ( .D(n8389), .CK(clk), .Q(reg_mem[1690]) );
  DFF_X1 reg_mem_reg_44__1_ ( .D(n8388), .CK(clk), .Q(reg_mem[1689]) );
  DFF_X1 reg_mem_reg_44__0_ ( .D(n8387), .CK(clk), .Q(reg_mem[1688]) );
  DFF_X1 reg_mem_reg_45__7_ ( .D(n7817), .CK(clk), .Q(reg_mem[1687]) );
  DFF_X1 reg_mem_reg_45__6_ ( .D(n7816), .CK(clk), .Q(reg_mem[1686]) );
  DFF_X1 reg_mem_reg_45__5_ ( .D(n7815), .CK(clk), .Q(reg_mem[1685]) );
  DFF_X1 reg_mem_reg_45__4_ ( .D(n7814), .CK(clk), .Q(reg_mem[1684]) );
  DFF_X1 reg_mem_reg_45__3_ ( .D(n7813), .CK(clk), .Q(reg_mem[1683]) );
  DFF_X1 reg_mem_reg_45__2_ ( .D(n7812), .CK(clk), .Q(reg_mem[1682]) );
  DFF_X1 reg_mem_reg_45__1_ ( .D(n7811), .CK(clk), .Q(reg_mem[1681]) );
  DFF_X1 reg_mem_reg_45__0_ ( .D(n7810), .CK(clk), .Q(reg_mem[1680]) );
  DFF_X1 reg_mem_reg_46__7_ ( .D(n8970), .CK(clk), .Q(reg_mem[1679]) );
  DFF_X1 reg_mem_reg_46__6_ ( .D(n8969), .CK(clk), .Q(reg_mem[1678]) );
  DFF_X1 reg_mem_reg_46__5_ ( .D(n8968), .CK(clk), .Q(reg_mem[1677]) );
  DFF_X1 reg_mem_reg_46__4_ ( .D(n8967), .CK(clk), .Q(reg_mem[1676]) );
  DFF_X1 reg_mem_reg_46__3_ ( .D(n8966), .CK(clk), .Q(reg_mem[1675]) );
  DFF_X1 reg_mem_reg_46__2_ ( .D(n8965), .CK(clk), .Q(reg_mem[1674]) );
  DFF_X1 reg_mem_reg_46__1_ ( .D(n8964), .CK(clk), .Q(reg_mem[1673]) );
  DFF_X1 reg_mem_reg_46__0_ ( .D(n8963), .CK(clk), .Q(reg_mem[1672]) );
  DFF_X1 reg_mem_reg_47__7_ ( .D(n7241), .CK(clk), .Q(reg_mem[1671]) );
  DFF_X1 reg_mem_reg_47__6_ ( .D(n7240), .CK(clk), .Q(reg_mem[1670]) );
  DFF_X1 reg_mem_reg_47__5_ ( .D(n7239), .CK(clk), .Q(reg_mem[1669]) );
  DFF_X1 reg_mem_reg_47__4_ ( .D(n7238), .CK(clk), .Q(reg_mem[1668]) );
  DFF_X1 reg_mem_reg_47__3_ ( .D(n7237), .CK(clk), .Q(reg_mem[1667]) );
  DFF_X1 reg_mem_reg_47__2_ ( .D(n7236), .CK(clk), .Q(reg_mem[1666]) );
  DFF_X1 reg_mem_reg_47__1_ ( .D(n7235), .CK(clk), .Q(reg_mem[1665]) );
  DFF_X1 reg_mem_reg_47__0_ ( .D(n7234), .CK(clk), .Q(reg_mem[1664]) );
  DFF_X1 reg_mem_reg_48__7_ ( .D(n7971), .CK(clk), .Q(reg_mem[1663]) );
  DFF_X1 reg_mem_reg_48__6_ ( .D(n7970), .CK(clk), .Q(reg_mem[1662]) );
  DFF_X1 reg_mem_reg_48__5_ ( .D(n7969), .CK(clk), .Q(reg_mem[1661]) );
  DFF_X1 reg_mem_reg_48__4_ ( .D(n7968), .CK(clk), .Q(reg_mem[1660]) );
  DFF_X1 reg_mem_reg_48__3_ ( .D(n7967), .CK(clk), .Q(reg_mem[1659]) );
  DFF_X1 reg_mem_reg_48__2_ ( .D(n7966), .CK(clk), .Q(reg_mem[1658]) );
  DFF_X1 reg_mem_reg_48__1_ ( .D(n7965), .CK(clk), .Q(reg_mem[1657]) );
  DFF_X1 reg_mem_reg_48__0_ ( .D(n7964), .CK(clk), .Q(reg_mem[1656]) );
  DFF_X1 reg_mem_reg_49__7_ ( .D(n7394), .CK(clk), .Q(reg_mem[1655]) );
  DFF_X1 reg_mem_reg_49__6_ ( .D(n7393), .CK(clk), .Q(reg_mem[1654]) );
  DFF_X1 reg_mem_reg_49__5_ ( .D(n7392), .CK(clk), .Q(reg_mem[1653]) );
  DFF_X1 reg_mem_reg_49__4_ ( .D(n7391), .CK(clk), .Q(reg_mem[1652]) );
  DFF_X1 reg_mem_reg_49__3_ ( .D(n7390), .CK(clk), .Q(reg_mem[1651]) );
  DFF_X1 reg_mem_reg_49__2_ ( .D(n7389), .CK(clk), .Q(reg_mem[1650]) );
  DFF_X1 reg_mem_reg_49__1_ ( .D(n7388), .CK(clk), .Q(reg_mem[1649]) );
  DFF_X1 reg_mem_reg_49__0_ ( .D(n7387), .CK(clk), .Q(reg_mem[1648]) );
  DFF_X1 reg_mem_reg_50__7_ ( .D(n8547), .CK(clk), .Q(reg_mem[1647]) );
  DFF_X1 reg_mem_reg_50__6_ ( .D(n8546), .CK(clk), .Q(reg_mem[1646]) );
  DFF_X1 reg_mem_reg_50__5_ ( .D(n8545), .CK(clk), .Q(reg_mem[1645]) );
  DFF_X1 reg_mem_reg_50__4_ ( .D(n8544), .CK(clk), .Q(reg_mem[1644]) );
  DFF_X1 reg_mem_reg_50__3_ ( .D(n8543), .CK(clk), .Q(reg_mem[1643]) );
  DFF_X1 reg_mem_reg_50__2_ ( .D(n8542), .CK(clk), .Q(reg_mem[1642]) );
  DFF_X1 reg_mem_reg_50__1_ ( .D(n8541), .CK(clk), .Q(reg_mem[1641]) );
  DFF_X1 reg_mem_reg_50__0_ ( .D(n8540), .CK(clk), .Q(reg_mem[1640]) );
  DFF_X1 reg_mem_reg_51__7_ ( .D(n6818), .CK(clk), .Q(reg_mem[1639]) );
  DFF_X1 reg_mem_reg_51__6_ ( .D(n6817), .CK(clk), .Q(reg_mem[1638]) );
  DFF_X1 reg_mem_reg_51__5_ ( .D(n6816), .CK(clk), .Q(reg_mem[1637]) );
  DFF_X1 reg_mem_reg_51__4_ ( .D(n6815), .CK(clk), .Q(reg_mem[1636]) );
  DFF_X1 reg_mem_reg_51__3_ ( .D(n6814), .CK(clk), .Q(reg_mem[1635]) );
  DFF_X1 reg_mem_reg_51__2_ ( .D(n6813), .CK(clk), .Q(reg_mem[1634]) );
  DFF_X1 reg_mem_reg_51__1_ ( .D(n6812), .CK(clk), .Q(reg_mem[1633]) );
  DFF_X1 reg_mem_reg_51__0_ ( .D(n6811), .CK(clk), .Q(reg_mem[1632]) );
  DFF_X1 reg_mem_reg_52__7_ ( .D(n8115), .CK(clk), .Q(reg_mem[1631]) );
  DFF_X1 reg_mem_reg_52__6_ ( .D(n8114), .CK(clk), .Q(reg_mem[1630]) );
  DFF_X1 reg_mem_reg_52__5_ ( .D(n8113), .CK(clk), .Q(reg_mem[1629]) );
  DFF_X1 reg_mem_reg_52__4_ ( .D(n8112), .CK(clk), .Q(reg_mem[1628]) );
  DFF_X1 reg_mem_reg_52__3_ ( .D(n8111), .CK(clk), .Q(reg_mem[1627]) );
  DFF_X1 reg_mem_reg_52__2_ ( .D(n8110), .CK(clk), .Q(reg_mem[1626]) );
  DFF_X1 reg_mem_reg_52__1_ ( .D(n8109), .CK(clk), .Q(reg_mem[1625]) );
  DFF_X1 reg_mem_reg_52__0_ ( .D(n8108), .CK(clk), .Q(reg_mem[1624]) );
  DFF_X1 reg_mem_reg_53__7_ ( .D(n7538), .CK(clk), .Q(reg_mem[1623]) );
  DFF_X1 reg_mem_reg_53__6_ ( .D(n7537), .CK(clk), .Q(reg_mem[1622]) );
  DFF_X1 reg_mem_reg_53__5_ ( .D(n7536), .CK(clk), .Q(reg_mem[1621]) );
  DFF_X1 reg_mem_reg_53__4_ ( .D(n7535), .CK(clk), .Q(reg_mem[1620]) );
  DFF_X1 reg_mem_reg_53__3_ ( .D(n7534), .CK(clk), .Q(reg_mem[1619]) );
  DFF_X1 reg_mem_reg_53__2_ ( .D(n7533), .CK(clk), .Q(reg_mem[1618]) );
  DFF_X1 reg_mem_reg_53__1_ ( .D(n7532), .CK(clk), .Q(reg_mem[1617]) );
  DFF_X1 reg_mem_reg_53__0_ ( .D(n7531), .CK(clk), .Q(reg_mem[1616]) );
  DFF_X1 reg_mem_reg_54__7_ ( .D(n8691), .CK(clk), .Q(reg_mem[1615]) );
  DFF_X1 reg_mem_reg_54__6_ ( .D(n8690), .CK(clk), .Q(reg_mem[1614]) );
  DFF_X1 reg_mem_reg_54__5_ ( .D(n8689), .CK(clk), .Q(reg_mem[1613]) );
  DFF_X1 reg_mem_reg_54__4_ ( .D(n8688), .CK(clk), .Q(reg_mem[1612]) );
  DFF_X1 reg_mem_reg_54__3_ ( .D(n8687), .CK(clk), .Q(reg_mem[1611]) );
  DFF_X1 reg_mem_reg_54__2_ ( .D(n8686), .CK(clk), .Q(reg_mem[1610]) );
  DFF_X1 reg_mem_reg_54__1_ ( .D(n8685), .CK(clk), .Q(reg_mem[1609]) );
  DFF_X1 reg_mem_reg_54__0_ ( .D(n8684), .CK(clk), .Q(reg_mem[1608]) );
  DFF_X1 reg_mem_reg_55__7_ ( .D(n6962), .CK(clk), .Q(reg_mem[1607]) );
  DFF_X1 reg_mem_reg_55__6_ ( .D(n6961), .CK(clk), .Q(reg_mem[1606]) );
  DFF_X1 reg_mem_reg_55__5_ ( .D(n6960), .CK(clk), .Q(reg_mem[1605]) );
  DFF_X1 reg_mem_reg_55__4_ ( .D(n6959), .CK(clk), .Q(reg_mem[1604]) );
  DFF_X1 reg_mem_reg_55__3_ ( .D(n6958), .CK(clk), .Q(reg_mem[1603]) );
  DFF_X1 reg_mem_reg_55__2_ ( .D(n6957), .CK(clk), .Q(reg_mem[1602]) );
  DFF_X1 reg_mem_reg_55__1_ ( .D(n6956), .CK(clk), .Q(reg_mem[1601]) );
  DFF_X1 reg_mem_reg_55__0_ ( .D(n6955), .CK(clk), .Q(reg_mem[1600]) );
  DFF_X1 reg_mem_reg_56__7_ ( .D(n8259), .CK(clk), .Q(reg_mem[1599]) );
  DFF_X1 reg_mem_reg_56__6_ ( .D(n8258), .CK(clk), .Q(reg_mem[1598]) );
  DFF_X1 reg_mem_reg_56__5_ ( .D(n8257), .CK(clk), .Q(reg_mem[1597]) );
  DFF_X1 reg_mem_reg_56__4_ ( .D(n8256), .CK(clk), .Q(reg_mem[1596]) );
  DFF_X1 reg_mem_reg_56__3_ ( .D(n8255), .CK(clk), .Q(reg_mem[1595]) );
  DFF_X1 reg_mem_reg_56__2_ ( .D(n8254), .CK(clk), .Q(reg_mem[1594]) );
  DFF_X1 reg_mem_reg_56__1_ ( .D(n8253), .CK(clk), .Q(reg_mem[1593]) );
  DFF_X1 reg_mem_reg_56__0_ ( .D(n8252), .CK(clk), .Q(reg_mem[1592]) );
  DFF_X1 reg_mem_reg_57__7_ ( .D(n7682), .CK(clk), .Q(reg_mem[1591]) );
  DFF_X1 reg_mem_reg_57__6_ ( .D(n7681), .CK(clk), .Q(reg_mem[1590]) );
  DFF_X1 reg_mem_reg_57__5_ ( .D(n7680), .CK(clk), .Q(reg_mem[1589]) );
  DFF_X1 reg_mem_reg_57__4_ ( .D(n7679), .CK(clk), .Q(reg_mem[1588]) );
  DFF_X1 reg_mem_reg_57__3_ ( .D(n7678), .CK(clk), .Q(reg_mem[1587]) );
  DFF_X1 reg_mem_reg_57__2_ ( .D(n7677), .CK(clk), .Q(reg_mem[1586]) );
  DFF_X1 reg_mem_reg_57__1_ ( .D(n7676), .CK(clk), .Q(reg_mem[1585]) );
  DFF_X1 reg_mem_reg_57__0_ ( .D(n7675), .CK(clk), .Q(reg_mem[1584]) );
  DFF_X1 reg_mem_reg_58__7_ ( .D(n8835), .CK(clk), .Q(reg_mem[1583]) );
  DFF_X1 reg_mem_reg_58__6_ ( .D(n8834), .CK(clk), .Q(reg_mem[1582]) );
  DFF_X1 reg_mem_reg_58__5_ ( .D(n8833), .CK(clk), .Q(reg_mem[1581]) );
  DFF_X1 reg_mem_reg_58__4_ ( .D(n8832), .CK(clk), .Q(reg_mem[1580]) );
  DFF_X1 reg_mem_reg_58__3_ ( .D(n8831), .CK(clk), .Q(reg_mem[1579]) );
  DFF_X1 reg_mem_reg_58__2_ ( .D(n8830), .CK(clk), .Q(reg_mem[1578]) );
  DFF_X1 reg_mem_reg_58__1_ ( .D(n8829), .CK(clk), .Q(reg_mem[1577]) );
  DFF_X1 reg_mem_reg_58__0_ ( .D(n8828), .CK(clk), .Q(reg_mem[1576]) );
  DFF_X1 reg_mem_reg_59__7_ ( .D(n7106), .CK(clk), .Q(reg_mem[1575]) );
  DFF_X1 reg_mem_reg_59__6_ ( .D(n7105), .CK(clk), .Q(reg_mem[1574]) );
  DFF_X1 reg_mem_reg_59__5_ ( .D(n7104), .CK(clk), .Q(reg_mem[1573]) );
  DFF_X1 reg_mem_reg_59__4_ ( .D(n7103), .CK(clk), .Q(reg_mem[1572]) );
  DFF_X1 reg_mem_reg_59__3_ ( .D(n7102), .CK(clk), .Q(reg_mem[1571]) );
  DFF_X1 reg_mem_reg_59__2_ ( .D(n7101), .CK(clk), .Q(reg_mem[1570]) );
  DFF_X1 reg_mem_reg_59__1_ ( .D(n7100), .CK(clk), .Q(reg_mem[1569]) );
  DFF_X1 reg_mem_reg_59__0_ ( .D(n7099), .CK(clk), .Q(reg_mem[1568]) );
  DFF_X1 reg_mem_reg_60__7_ ( .D(n8403), .CK(clk), .Q(reg_mem[1567]) );
  DFF_X1 reg_mem_reg_60__6_ ( .D(n8402), .CK(clk), .Q(reg_mem[1566]) );
  DFF_X1 reg_mem_reg_60__5_ ( .D(n8401), .CK(clk), .Q(reg_mem[1565]) );
  DFF_X1 reg_mem_reg_60__4_ ( .D(n8400), .CK(clk), .Q(reg_mem[1564]) );
  DFF_X1 reg_mem_reg_60__3_ ( .D(n8399), .CK(clk), .Q(reg_mem[1563]) );
  DFF_X1 reg_mem_reg_60__2_ ( .D(n8398), .CK(clk), .Q(reg_mem[1562]) );
  DFF_X1 reg_mem_reg_60__1_ ( .D(n8397), .CK(clk), .Q(reg_mem[1561]) );
  DFF_X1 reg_mem_reg_60__0_ ( .D(n8396), .CK(clk), .Q(reg_mem[1560]) );
  DFF_X1 reg_mem_reg_61__7_ ( .D(n7826), .CK(clk), .Q(reg_mem[1559]) );
  DFF_X1 reg_mem_reg_61__6_ ( .D(n7825), .CK(clk), .Q(reg_mem[1558]) );
  DFF_X1 reg_mem_reg_61__5_ ( .D(n7824), .CK(clk), .Q(reg_mem[1557]) );
  DFF_X1 reg_mem_reg_61__4_ ( .D(n7823), .CK(clk), .Q(reg_mem[1556]) );
  DFF_X1 reg_mem_reg_61__3_ ( .D(n7822), .CK(clk), .Q(reg_mem[1555]) );
  DFF_X1 reg_mem_reg_61__2_ ( .D(n7821), .CK(clk), .Q(reg_mem[1554]) );
  DFF_X1 reg_mem_reg_61__1_ ( .D(n7820), .CK(clk), .Q(reg_mem[1553]) );
  DFF_X1 reg_mem_reg_61__0_ ( .D(n7819), .CK(clk), .Q(reg_mem[1552]) );
  DFF_X1 reg_mem_reg_62__7_ ( .D(n8979), .CK(clk), .Q(reg_mem[1551]) );
  DFF_X1 reg_mem_reg_62__6_ ( .D(n8978), .CK(clk), .Q(reg_mem[1550]) );
  DFF_X1 reg_mem_reg_62__5_ ( .D(n8977), .CK(clk), .Q(reg_mem[1549]) );
  DFF_X1 reg_mem_reg_62__4_ ( .D(n8976), .CK(clk), .Q(reg_mem[1548]) );
  DFF_X1 reg_mem_reg_62__3_ ( .D(n8975), .CK(clk), .Q(reg_mem[1547]) );
  DFF_X1 reg_mem_reg_62__2_ ( .D(n8974), .CK(clk), .Q(reg_mem[1546]) );
  DFF_X1 reg_mem_reg_62__1_ ( .D(n8973), .CK(clk), .Q(reg_mem[1545]) );
  DFF_X1 reg_mem_reg_62__0_ ( .D(n8972), .CK(clk), .Q(reg_mem[1544]) );
  DFF_X1 reg_mem_reg_63__7_ ( .D(n7250), .CK(clk), .Q(reg_mem[1543]) );
  DFF_X1 reg_mem_reg_63__6_ ( .D(n7249), .CK(clk), .Q(reg_mem[1542]) );
  DFF_X1 reg_mem_reg_63__5_ ( .D(n7248), .CK(clk), .Q(reg_mem[1541]) );
  DFF_X1 reg_mem_reg_63__4_ ( .D(n7247), .CK(clk), .Q(reg_mem[1540]) );
  DFF_X1 reg_mem_reg_63__3_ ( .D(n7246), .CK(clk), .Q(reg_mem[1539]) );
  DFF_X1 reg_mem_reg_63__2_ ( .D(n7245), .CK(clk), .Q(reg_mem[1538]) );
  DFF_X1 reg_mem_reg_63__1_ ( .D(n7244), .CK(clk), .Q(reg_mem[1537]) );
  DFF_X1 reg_mem_reg_63__0_ ( .D(n7243), .CK(clk), .Q(reg_mem[1536]) );
  DFF_X1 reg_mem_reg_64__7_ ( .D(n7980), .CK(clk), .Q(reg_mem[1535]) );
  DFF_X1 reg_mem_reg_64__6_ ( .D(n7979), .CK(clk), .Q(reg_mem[1534]) );
  DFF_X1 reg_mem_reg_64__5_ ( .D(n7978), .CK(clk), .Q(reg_mem[1533]) );
  DFF_X1 reg_mem_reg_64__4_ ( .D(n7977), .CK(clk), .Q(reg_mem[1532]) );
  DFF_X1 reg_mem_reg_64__3_ ( .D(n7976), .CK(clk), .Q(reg_mem[1531]) );
  DFF_X1 reg_mem_reg_64__2_ ( .D(n7975), .CK(clk), .Q(reg_mem[1530]) );
  DFF_X1 reg_mem_reg_64__1_ ( .D(n7974), .CK(clk), .Q(reg_mem[1529]) );
  DFF_X1 reg_mem_reg_64__0_ ( .D(n7973), .CK(clk), .Q(reg_mem[1528]) );
  DFF_X1 reg_mem_reg_65__7_ ( .D(n7403), .CK(clk), .Q(reg_mem[1527]) );
  DFF_X1 reg_mem_reg_65__6_ ( .D(n7402), .CK(clk), .Q(reg_mem[1526]) );
  DFF_X1 reg_mem_reg_65__5_ ( .D(n7401), .CK(clk), .Q(reg_mem[1525]) );
  DFF_X1 reg_mem_reg_65__4_ ( .D(n7400), .CK(clk), .Q(reg_mem[1524]) );
  DFF_X1 reg_mem_reg_65__3_ ( .D(n7399), .CK(clk), .Q(reg_mem[1523]) );
  DFF_X1 reg_mem_reg_65__2_ ( .D(n7398), .CK(clk), .Q(reg_mem[1522]) );
  DFF_X1 reg_mem_reg_65__1_ ( .D(n7397), .CK(clk), .Q(reg_mem[1521]) );
  DFF_X1 reg_mem_reg_65__0_ ( .D(n7396), .CK(clk), .Q(reg_mem[1520]) );
  DFF_X1 reg_mem_reg_66__7_ ( .D(n8556), .CK(clk), .Q(reg_mem[1519]) );
  DFF_X1 reg_mem_reg_66__6_ ( .D(n8555), .CK(clk), .Q(reg_mem[1518]) );
  DFF_X1 reg_mem_reg_66__5_ ( .D(n8554), .CK(clk), .Q(reg_mem[1517]) );
  DFF_X1 reg_mem_reg_66__4_ ( .D(n8553), .CK(clk), .Q(reg_mem[1516]) );
  DFF_X1 reg_mem_reg_66__3_ ( .D(n8552), .CK(clk), .Q(reg_mem[1515]) );
  DFF_X1 reg_mem_reg_66__2_ ( .D(n8551), .CK(clk), .Q(reg_mem[1514]) );
  DFF_X1 reg_mem_reg_66__1_ ( .D(n8550), .CK(clk), .Q(reg_mem[1513]) );
  DFF_X1 reg_mem_reg_66__0_ ( .D(n8549), .CK(clk), .Q(reg_mem[1512]) );
  DFF_X1 reg_mem_reg_67__7_ ( .D(n6827), .CK(clk), .Q(reg_mem[1511]) );
  DFF_X1 reg_mem_reg_67__6_ ( .D(n6826), .CK(clk), .Q(reg_mem[1510]) );
  DFF_X1 reg_mem_reg_67__5_ ( .D(n6825), .CK(clk), .Q(reg_mem[1509]) );
  DFF_X1 reg_mem_reg_67__4_ ( .D(n6824), .CK(clk), .Q(reg_mem[1508]) );
  DFF_X1 reg_mem_reg_67__3_ ( .D(n6823), .CK(clk), .Q(reg_mem[1507]) );
  DFF_X1 reg_mem_reg_67__2_ ( .D(n6822), .CK(clk), .Q(reg_mem[1506]) );
  DFF_X1 reg_mem_reg_67__1_ ( .D(n6821), .CK(clk), .Q(reg_mem[1505]) );
  DFF_X1 reg_mem_reg_67__0_ ( .D(n6820), .CK(clk), .Q(reg_mem[1504]) );
  DFF_X1 reg_mem_reg_68__7_ ( .D(n8124), .CK(clk), .Q(reg_mem[1503]) );
  DFF_X1 reg_mem_reg_68__6_ ( .D(n8123), .CK(clk), .Q(reg_mem[1502]) );
  DFF_X1 reg_mem_reg_68__5_ ( .D(n8122), .CK(clk), .Q(reg_mem[1501]) );
  DFF_X1 reg_mem_reg_68__4_ ( .D(n8121), .CK(clk), .Q(reg_mem[1500]) );
  DFF_X1 reg_mem_reg_68__3_ ( .D(n8120), .CK(clk), .Q(reg_mem[1499]) );
  DFF_X1 reg_mem_reg_68__2_ ( .D(n8119), .CK(clk), .Q(reg_mem[1498]) );
  DFF_X1 reg_mem_reg_68__1_ ( .D(n8118), .CK(clk), .Q(reg_mem[1497]) );
  DFF_X1 reg_mem_reg_68__0_ ( .D(n8117), .CK(clk), .Q(reg_mem[1496]) );
  DFF_X1 reg_mem_reg_69__7_ ( .D(n7547), .CK(clk), .Q(reg_mem[1495]) );
  DFF_X1 reg_mem_reg_69__6_ ( .D(n7546), .CK(clk), .Q(reg_mem[1494]) );
  DFF_X1 reg_mem_reg_69__5_ ( .D(n7545), .CK(clk), .Q(reg_mem[1493]) );
  DFF_X1 reg_mem_reg_69__4_ ( .D(n7544), .CK(clk), .Q(reg_mem[1492]) );
  DFF_X1 reg_mem_reg_69__3_ ( .D(n7543), .CK(clk), .Q(reg_mem[1491]) );
  DFF_X1 reg_mem_reg_69__2_ ( .D(n7542), .CK(clk), .Q(reg_mem[1490]) );
  DFF_X1 reg_mem_reg_69__1_ ( .D(n7541), .CK(clk), .Q(reg_mem[1489]) );
  DFF_X1 reg_mem_reg_69__0_ ( .D(n7540), .CK(clk), .Q(reg_mem[1488]) );
  DFF_X1 reg_mem_reg_70__7_ ( .D(n8700), .CK(clk), .Q(reg_mem[1487]) );
  DFF_X1 reg_mem_reg_70__6_ ( .D(n8699), .CK(clk), .Q(reg_mem[1486]) );
  DFF_X1 reg_mem_reg_70__5_ ( .D(n8698), .CK(clk), .Q(reg_mem[1485]) );
  DFF_X1 reg_mem_reg_70__4_ ( .D(n8697), .CK(clk), .Q(reg_mem[1484]) );
  DFF_X1 reg_mem_reg_70__3_ ( .D(n8696), .CK(clk), .Q(reg_mem[1483]) );
  DFF_X1 reg_mem_reg_70__2_ ( .D(n8695), .CK(clk), .Q(reg_mem[1482]) );
  DFF_X1 reg_mem_reg_70__1_ ( .D(n8694), .CK(clk), .Q(reg_mem[1481]) );
  DFF_X1 reg_mem_reg_70__0_ ( .D(n8693), .CK(clk), .Q(reg_mem[1480]) );
  DFF_X1 reg_mem_reg_71__7_ ( .D(n6971), .CK(clk), .Q(reg_mem[1479]) );
  DFF_X1 reg_mem_reg_71__6_ ( .D(n6970), .CK(clk), .Q(reg_mem[1478]) );
  DFF_X1 reg_mem_reg_71__5_ ( .D(n6969), .CK(clk), .Q(reg_mem[1477]) );
  DFF_X1 reg_mem_reg_71__4_ ( .D(n6968), .CK(clk), .Q(reg_mem[1476]) );
  DFF_X1 reg_mem_reg_71__3_ ( .D(n6967), .CK(clk), .Q(reg_mem[1475]) );
  DFF_X1 reg_mem_reg_71__2_ ( .D(n6966), .CK(clk), .Q(reg_mem[1474]) );
  DFF_X1 reg_mem_reg_71__1_ ( .D(n6965), .CK(clk), .Q(reg_mem[1473]) );
  DFF_X1 reg_mem_reg_71__0_ ( .D(n6964), .CK(clk), .Q(reg_mem[1472]) );
  DFF_X1 reg_mem_reg_72__7_ ( .D(n8268), .CK(clk), .Q(reg_mem[1471]) );
  DFF_X1 reg_mem_reg_72__6_ ( .D(n8267), .CK(clk), .Q(reg_mem[1470]) );
  DFF_X1 reg_mem_reg_72__5_ ( .D(n8266), .CK(clk), .Q(reg_mem[1469]) );
  DFF_X1 reg_mem_reg_72__4_ ( .D(n8265), .CK(clk), .Q(reg_mem[1468]) );
  DFF_X1 reg_mem_reg_72__3_ ( .D(n8264), .CK(clk), .Q(reg_mem[1467]) );
  DFF_X1 reg_mem_reg_72__2_ ( .D(n8263), .CK(clk), .Q(reg_mem[1466]) );
  DFF_X1 reg_mem_reg_72__1_ ( .D(n8262), .CK(clk), .Q(reg_mem[1465]) );
  DFF_X1 reg_mem_reg_72__0_ ( .D(n8261), .CK(clk), .Q(reg_mem[1464]) );
  DFF_X1 reg_mem_reg_73__7_ ( .D(n7691), .CK(clk), .Q(reg_mem[1463]) );
  DFF_X1 reg_mem_reg_73__6_ ( .D(n7690), .CK(clk), .Q(reg_mem[1462]) );
  DFF_X1 reg_mem_reg_73__5_ ( .D(n7689), .CK(clk), .Q(reg_mem[1461]) );
  DFF_X1 reg_mem_reg_73__4_ ( .D(n7688), .CK(clk), .Q(reg_mem[1460]) );
  DFF_X1 reg_mem_reg_73__3_ ( .D(n7687), .CK(clk), .Q(reg_mem[1459]) );
  DFF_X1 reg_mem_reg_73__2_ ( .D(n7686), .CK(clk), .Q(reg_mem[1458]) );
  DFF_X1 reg_mem_reg_73__1_ ( .D(n7685), .CK(clk), .Q(reg_mem[1457]) );
  DFF_X1 reg_mem_reg_73__0_ ( .D(n7684), .CK(clk), .Q(reg_mem[1456]) );
  DFF_X1 reg_mem_reg_74__7_ ( .D(n8844), .CK(clk), .Q(reg_mem[1455]) );
  DFF_X1 reg_mem_reg_74__6_ ( .D(n8843), .CK(clk), .Q(reg_mem[1454]) );
  DFF_X1 reg_mem_reg_74__5_ ( .D(n8842), .CK(clk), .Q(reg_mem[1453]) );
  DFF_X1 reg_mem_reg_74__4_ ( .D(n8841), .CK(clk), .Q(reg_mem[1452]) );
  DFF_X1 reg_mem_reg_74__3_ ( .D(n8840), .CK(clk), .Q(reg_mem[1451]) );
  DFF_X1 reg_mem_reg_74__2_ ( .D(n8839), .CK(clk), .Q(reg_mem[1450]) );
  DFF_X1 reg_mem_reg_74__1_ ( .D(n8838), .CK(clk), .Q(reg_mem[1449]) );
  DFF_X1 reg_mem_reg_74__0_ ( .D(n8837), .CK(clk), .Q(reg_mem[1448]) );
  DFF_X1 reg_mem_reg_75__7_ ( .D(n7115), .CK(clk), .Q(reg_mem[1447]) );
  DFF_X1 reg_mem_reg_75__6_ ( .D(n7114), .CK(clk), .Q(reg_mem[1446]) );
  DFF_X1 reg_mem_reg_75__5_ ( .D(n7113), .CK(clk), .Q(reg_mem[1445]) );
  DFF_X1 reg_mem_reg_75__4_ ( .D(n7112), .CK(clk), .Q(reg_mem[1444]) );
  DFF_X1 reg_mem_reg_75__3_ ( .D(n7111), .CK(clk), .Q(reg_mem[1443]) );
  DFF_X1 reg_mem_reg_75__2_ ( .D(n7110), .CK(clk), .Q(reg_mem[1442]) );
  DFF_X1 reg_mem_reg_75__1_ ( .D(n7109), .CK(clk), .Q(reg_mem[1441]) );
  DFF_X1 reg_mem_reg_75__0_ ( .D(n7108), .CK(clk), .Q(reg_mem[1440]) );
  DFF_X1 reg_mem_reg_76__7_ ( .D(n8412), .CK(clk), .Q(reg_mem[1439]) );
  DFF_X1 reg_mem_reg_76__6_ ( .D(n8411), .CK(clk), .Q(reg_mem[1438]) );
  DFF_X1 reg_mem_reg_76__5_ ( .D(n8410), .CK(clk), .Q(reg_mem[1437]) );
  DFF_X1 reg_mem_reg_76__4_ ( .D(n8409), .CK(clk), .Q(reg_mem[1436]) );
  DFF_X1 reg_mem_reg_76__3_ ( .D(n8408), .CK(clk), .Q(reg_mem[1435]) );
  DFF_X1 reg_mem_reg_76__2_ ( .D(n8407), .CK(clk), .Q(reg_mem[1434]) );
  DFF_X1 reg_mem_reg_76__1_ ( .D(n8406), .CK(clk), .Q(reg_mem[1433]) );
  DFF_X1 reg_mem_reg_76__0_ ( .D(n8405), .CK(clk), .Q(reg_mem[1432]) );
  DFF_X1 reg_mem_reg_77__7_ ( .D(n7835), .CK(clk), .Q(reg_mem[1431]) );
  DFF_X1 reg_mem_reg_77__6_ ( .D(n7834), .CK(clk), .Q(reg_mem[1430]) );
  DFF_X1 reg_mem_reg_77__5_ ( .D(n7833), .CK(clk), .Q(reg_mem[1429]) );
  DFF_X1 reg_mem_reg_77__4_ ( .D(n7832), .CK(clk), .Q(reg_mem[1428]) );
  DFF_X1 reg_mem_reg_77__3_ ( .D(n7831), .CK(clk), .Q(reg_mem[1427]) );
  DFF_X1 reg_mem_reg_77__2_ ( .D(n7830), .CK(clk), .Q(reg_mem[1426]) );
  DFF_X1 reg_mem_reg_77__1_ ( .D(n7829), .CK(clk), .Q(reg_mem[1425]) );
  DFF_X1 reg_mem_reg_77__0_ ( .D(n7828), .CK(clk), .Q(reg_mem[1424]) );
  DFF_X1 reg_mem_reg_78__7_ ( .D(n8988), .CK(clk), .Q(reg_mem[1423]) );
  DFF_X1 reg_mem_reg_78__6_ ( .D(n8987), .CK(clk), .Q(reg_mem[1422]) );
  DFF_X1 reg_mem_reg_78__5_ ( .D(n8986), .CK(clk), .Q(reg_mem[1421]) );
  DFF_X1 reg_mem_reg_78__4_ ( .D(n8985), .CK(clk), .Q(reg_mem[1420]) );
  DFF_X1 reg_mem_reg_78__3_ ( .D(n8984), .CK(clk), .Q(reg_mem[1419]) );
  DFF_X1 reg_mem_reg_78__2_ ( .D(n8983), .CK(clk), .Q(reg_mem[1418]) );
  DFF_X1 reg_mem_reg_78__1_ ( .D(n8982), .CK(clk), .Q(reg_mem[1417]) );
  DFF_X1 reg_mem_reg_78__0_ ( .D(n8981), .CK(clk), .Q(reg_mem[1416]) );
  DFF_X1 reg_mem_reg_79__7_ ( .D(n7259), .CK(clk), .Q(reg_mem[1415]) );
  DFF_X1 reg_mem_reg_79__6_ ( .D(n7258), .CK(clk), .Q(reg_mem[1414]) );
  DFF_X1 reg_mem_reg_79__5_ ( .D(n7257), .CK(clk), .Q(reg_mem[1413]) );
  DFF_X1 reg_mem_reg_79__4_ ( .D(n7256), .CK(clk), .Q(reg_mem[1412]) );
  DFF_X1 reg_mem_reg_79__3_ ( .D(n7255), .CK(clk), .Q(reg_mem[1411]) );
  DFF_X1 reg_mem_reg_79__2_ ( .D(n7254), .CK(clk), .Q(reg_mem[1410]) );
  DFF_X1 reg_mem_reg_79__1_ ( .D(n7253), .CK(clk), .Q(reg_mem[1409]) );
  DFF_X1 reg_mem_reg_79__0_ ( .D(n7252), .CK(clk), .Q(reg_mem[1408]) );
  DFF_X1 reg_mem_reg_80__7_ ( .D(n7989), .CK(clk), .Q(reg_mem[1407]) );
  DFF_X1 reg_mem_reg_80__6_ ( .D(n7988), .CK(clk), .Q(reg_mem[1406]) );
  DFF_X1 reg_mem_reg_80__5_ ( .D(n7987), .CK(clk), .Q(reg_mem[1405]) );
  DFF_X1 reg_mem_reg_80__4_ ( .D(n7986), .CK(clk), .Q(reg_mem[1404]) );
  DFF_X1 reg_mem_reg_80__3_ ( .D(n7985), .CK(clk), .Q(reg_mem[1403]) );
  DFF_X1 reg_mem_reg_80__2_ ( .D(n7984), .CK(clk), .Q(reg_mem[1402]) );
  DFF_X1 reg_mem_reg_80__1_ ( .D(n7983), .CK(clk), .Q(reg_mem[1401]) );
  DFF_X1 reg_mem_reg_80__0_ ( .D(n7982), .CK(clk), .Q(reg_mem[1400]) );
  DFF_X1 reg_mem_reg_81__7_ ( .D(n7412), .CK(clk), .Q(reg_mem[1399]) );
  DFF_X1 reg_mem_reg_81__6_ ( .D(n7411), .CK(clk), .Q(reg_mem[1398]) );
  DFF_X1 reg_mem_reg_81__5_ ( .D(n7410), .CK(clk), .Q(reg_mem[1397]) );
  DFF_X1 reg_mem_reg_81__4_ ( .D(n7409), .CK(clk), .Q(reg_mem[1396]) );
  DFF_X1 reg_mem_reg_81__3_ ( .D(n7408), .CK(clk), .Q(reg_mem[1395]) );
  DFF_X1 reg_mem_reg_81__2_ ( .D(n7407), .CK(clk), .Q(reg_mem[1394]) );
  DFF_X1 reg_mem_reg_81__1_ ( .D(n7406), .CK(clk), .Q(reg_mem[1393]) );
  DFF_X1 reg_mem_reg_81__0_ ( .D(n7405), .CK(clk), .Q(reg_mem[1392]) );
  DFF_X1 reg_mem_reg_82__7_ ( .D(n8565), .CK(clk), .Q(reg_mem[1391]) );
  DFF_X1 reg_mem_reg_82__6_ ( .D(n8564), .CK(clk), .Q(reg_mem[1390]) );
  DFF_X1 reg_mem_reg_82__5_ ( .D(n8563), .CK(clk), .Q(reg_mem[1389]) );
  DFF_X1 reg_mem_reg_82__4_ ( .D(n8562), .CK(clk), .Q(reg_mem[1388]) );
  DFF_X1 reg_mem_reg_82__3_ ( .D(n8561), .CK(clk), .Q(reg_mem[1387]) );
  DFF_X1 reg_mem_reg_82__2_ ( .D(n8560), .CK(clk), .Q(reg_mem[1386]) );
  DFF_X1 reg_mem_reg_82__1_ ( .D(n8559), .CK(clk), .Q(reg_mem[1385]) );
  DFF_X1 reg_mem_reg_82__0_ ( .D(n8558), .CK(clk), .Q(reg_mem[1384]) );
  DFF_X1 reg_mem_reg_83__7_ ( .D(n6836), .CK(clk), .Q(reg_mem[1383]) );
  DFF_X1 reg_mem_reg_83__6_ ( .D(n6835), .CK(clk), .Q(reg_mem[1382]) );
  DFF_X1 reg_mem_reg_83__5_ ( .D(n6834), .CK(clk), .Q(reg_mem[1381]) );
  DFF_X1 reg_mem_reg_83__4_ ( .D(n6833), .CK(clk), .Q(reg_mem[1380]) );
  DFF_X1 reg_mem_reg_83__3_ ( .D(n6832), .CK(clk), .Q(reg_mem[1379]) );
  DFF_X1 reg_mem_reg_83__2_ ( .D(n6831), .CK(clk), .Q(reg_mem[1378]) );
  DFF_X1 reg_mem_reg_83__1_ ( .D(n6830), .CK(clk), .Q(reg_mem[1377]) );
  DFF_X1 reg_mem_reg_83__0_ ( .D(n6829), .CK(clk), .Q(reg_mem[1376]) );
  DFF_X1 reg_mem_reg_84__7_ ( .D(n8133), .CK(clk), .Q(reg_mem[1375]) );
  DFF_X1 reg_mem_reg_84__6_ ( .D(n8132), .CK(clk), .Q(reg_mem[1374]) );
  DFF_X1 reg_mem_reg_84__5_ ( .D(n8131), .CK(clk), .Q(reg_mem[1373]) );
  DFF_X1 reg_mem_reg_84__4_ ( .D(n8130), .CK(clk), .Q(reg_mem[1372]) );
  DFF_X1 reg_mem_reg_84__3_ ( .D(n8129), .CK(clk), .Q(reg_mem[1371]) );
  DFF_X1 reg_mem_reg_84__2_ ( .D(n8128), .CK(clk), .Q(reg_mem[1370]) );
  DFF_X1 reg_mem_reg_84__1_ ( .D(n8127), .CK(clk), .Q(reg_mem[1369]) );
  DFF_X1 reg_mem_reg_84__0_ ( .D(n8126), .CK(clk), .Q(reg_mem[1368]) );
  DFF_X1 reg_mem_reg_85__7_ ( .D(n7556), .CK(clk), .Q(reg_mem[1367]) );
  DFF_X1 reg_mem_reg_85__6_ ( .D(n7555), .CK(clk), .Q(reg_mem[1366]) );
  DFF_X1 reg_mem_reg_85__5_ ( .D(n7554), .CK(clk), .Q(reg_mem[1365]) );
  DFF_X1 reg_mem_reg_85__4_ ( .D(n7553), .CK(clk), .Q(reg_mem[1364]) );
  DFF_X1 reg_mem_reg_85__3_ ( .D(n7552), .CK(clk), .Q(reg_mem[1363]) );
  DFF_X1 reg_mem_reg_85__2_ ( .D(n7551), .CK(clk), .Q(reg_mem[1362]) );
  DFF_X1 reg_mem_reg_85__1_ ( .D(n7550), .CK(clk), .Q(reg_mem[1361]) );
  DFF_X1 reg_mem_reg_85__0_ ( .D(n7549), .CK(clk), .Q(reg_mem[1360]) );
  DFF_X1 reg_mem_reg_86__7_ ( .D(n8709), .CK(clk), .Q(reg_mem[1359]) );
  DFF_X1 reg_mem_reg_86__6_ ( .D(n8708), .CK(clk), .Q(reg_mem[1358]) );
  DFF_X1 reg_mem_reg_86__5_ ( .D(n8707), .CK(clk), .Q(reg_mem[1357]) );
  DFF_X1 reg_mem_reg_86__4_ ( .D(n8706), .CK(clk), .Q(reg_mem[1356]) );
  DFF_X1 reg_mem_reg_86__3_ ( .D(n8705), .CK(clk), .Q(reg_mem[1355]) );
  DFF_X1 reg_mem_reg_86__2_ ( .D(n8704), .CK(clk), .Q(reg_mem[1354]) );
  DFF_X1 reg_mem_reg_86__1_ ( .D(n8703), .CK(clk), .Q(reg_mem[1353]) );
  DFF_X1 reg_mem_reg_86__0_ ( .D(n8702), .CK(clk), .Q(reg_mem[1352]) );
  DFF_X1 reg_mem_reg_87__7_ ( .D(n6980), .CK(clk), .Q(reg_mem[1351]) );
  DFF_X1 reg_mem_reg_87__6_ ( .D(n6979), .CK(clk), .Q(reg_mem[1350]) );
  DFF_X1 reg_mem_reg_87__5_ ( .D(n6978), .CK(clk), .Q(reg_mem[1349]) );
  DFF_X1 reg_mem_reg_87__4_ ( .D(n6977), .CK(clk), .Q(reg_mem[1348]) );
  DFF_X1 reg_mem_reg_87__3_ ( .D(n6976), .CK(clk), .Q(reg_mem[1347]) );
  DFF_X1 reg_mem_reg_87__2_ ( .D(n6975), .CK(clk), .Q(reg_mem[1346]) );
  DFF_X1 reg_mem_reg_87__1_ ( .D(n6974), .CK(clk), .Q(reg_mem[1345]) );
  DFF_X1 reg_mem_reg_87__0_ ( .D(n6973), .CK(clk), .Q(reg_mem[1344]) );
  DFF_X1 reg_mem_reg_88__7_ ( .D(n8277), .CK(clk), .Q(reg_mem[1343]) );
  DFF_X1 reg_mem_reg_88__6_ ( .D(n8276), .CK(clk), .Q(reg_mem[1342]) );
  DFF_X1 reg_mem_reg_88__5_ ( .D(n8275), .CK(clk), .Q(reg_mem[1341]) );
  DFF_X1 reg_mem_reg_88__4_ ( .D(n8274), .CK(clk), .Q(reg_mem[1340]) );
  DFF_X1 reg_mem_reg_88__3_ ( .D(n8273), .CK(clk), .Q(reg_mem[1339]) );
  DFF_X1 reg_mem_reg_88__2_ ( .D(n8272), .CK(clk), .Q(reg_mem[1338]) );
  DFF_X1 reg_mem_reg_88__1_ ( .D(n8271), .CK(clk), .Q(reg_mem[1337]) );
  DFF_X1 reg_mem_reg_88__0_ ( .D(n8270), .CK(clk), .Q(reg_mem[1336]) );
  DFF_X1 reg_mem_reg_89__7_ ( .D(n7700), .CK(clk), .Q(reg_mem[1335]) );
  DFF_X1 reg_mem_reg_89__6_ ( .D(n7699), .CK(clk), .Q(reg_mem[1334]) );
  DFF_X1 reg_mem_reg_89__5_ ( .D(n7698), .CK(clk), .Q(reg_mem[1333]) );
  DFF_X1 reg_mem_reg_89__4_ ( .D(n7697), .CK(clk), .Q(reg_mem[1332]) );
  DFF_X1 reg_mem_reg_89__3_ ( .D(n7696), .CK(clk), .Q(reg_mem[1331]) );
  DFF_X1 reg_mem_reg_89__2_ ( .D(n7695), .CK(clk), .Q(reg_mem[1330]) );
  DFF_X1 reg_mem_reg_89__1_ ( .D(n7694), .CK(clk), .Q(reg_mem[1329]) );
  DFF_X1 reg_mem_reg_89__0_ ( .D(n7693), .CK(clk), .Q(reg_mem[1328]) );
  DFF_X1 reg_mem_reg_90__7_ ( .D(n8853), .CK(clk), .Q(reg_mem[1327]) );
  DFF_X1 reg_mem_reg_90__6_ ( .D(n8852), .CK(clk), .Q(reg_mem[1326]) );
  DFF_X1 reg_mem_reg_90__5_ ( .D(n8851), .CK(clk), .Q(reg_mem[1325]) );
  DFF_X1 reg_mem_reg_90__4_ ( .D(n8850), .CK(clk), .Q(reg_mem[1324]) );
  DFF_X1 reg_mem_reg_90__3_ ( .D(n8849), .CK(clk), .Q(reg_mem[1323]) );
  DFF_X1 reg_mem_reg_90__2_ ( .D(n8848), .CK(clk), .Q(reg_mem[1322]) );
  DFF_X1 reg_mem_reg_90__1_ ( .D(n8847), .CK(clk), .Q(reg_mem[1321]) );
  DFF_X1 reg_mem_reg_90__0_ ( .D(n8846), .CK(clk), .Q(reg_mem[1320]) );
  DFF_X1 reg_mem_reg_91__7_ ( .D(n7124), .CK(clk), .Q(reg_mem[1319]) );
  DFF_X1 reg_mem_reg_91__6_ ( .D(n7123), .CK(clk), .Q(reg_mem[1318]) );
  DFF_X1 reg_mem_reg_91__5_ ( .D(n7122), .CK(clk), .Q(reg_mem[1317]) );
  DFF_X1 reg_mem_reg_91__4_ ( .D(n7121), .CK(clk), .Q(reg_mem[1316]) );
  DFF_X1 reg_mem_reg_91__3_ ( .D(n7120), .CK(clk), .Q(reg_mem[1315]) );
  DFF_X1 reg_mem_reg_91__2_ ( .D(n7119), .CK(clk), .Q(reg_mem[1314]) );
  DFF_X1 reg_mem_reg_91__1_ ( .D(n7118), .CK(clk), .Q(reg_mem[1313]) );
  DFF_X1 reg_mem_reg_91__0_ ( .D(n7117), .CK(clk), .Q(reg_mem[1312]) );
  DFF_X1 reg_mem_reg_92__7_ ( .D(n8421), .CK(clk), .Q(reg_mem[1311]) );
  DFF_X1 reg_mem_reg_92__6_ ( .D(n8420), .CK(clk), .Q(reg_mem[1310]) );
  DFF_X1 reg_mem_reg_92__5_ ( .D(n8419), .CK(clk), .Q(reg_mem[1309]) );
  DFF_X1 reg_mem_reg_92__4_ ( .D(n8418), .CK(clk), .Q(reg_mem[1308]) );
  DFF_X1 reg_mem_reg_92__3_ ( .D(n8417), .CK(clk), .Q(reg_mem[1307]) );
  DFF_X1 reg_mem_reg_92__2_ ( .D(n8416), .CK(clk), .Q(reg_mem[1306]) );
  DFF_X1 reg_mem_reg_92__1_ ( .D(n8415), .CK(clk), .Q(reg_mem[1305]) );
  DFF_X1 reg_mem_reg_92__0_ ( .D(n8414), .CK(clk), .Q(reg_mem[1304]) );
  DFF_X1 reg_mem_reg_93__7_ ( .D(n7844), .CK(clk), .Q(reg_mem[1303]) );
  DFF_X1 reg_mem_reg_93__6_ ( .D(n7843), .CK(clk), .Q(reg_mem[1302]) );
  DFF_X1 reg_mem_reg_93__5_ ( .D(n7842), .CK(clk), .Q(reg_mem[1301]) );
  DFF_X1 reg_mem_reg_93__4_ ( .D(n7841), .CK(clk), .Q(reg_mem[1300]) );
  DFF_X1 reg_mem_reg_93__3_ ( .D(n7840), .CK(clk), .Q(reg_mem[1299]) );
  DFF_X1 reg_mem_reg_93__2_ ( .D(n7839), .CK(clk), .Q(reg_mem[1298]) );
  DFF_X1 reg_mem_reg_93__1_ ( .D(n7838), .CK(clk), .Q(reg_mem[1297]) );
  DFF_X1 reg_mem_reg_93__0_ ( .D(n7837), .CK(clk), .Q(reg_mem[1296]) );
  DFF_X1 reg_mem_reg_94__7_ ( .D(n8997), .CK(clk), .Q(reg_mem[1295]) );
  DFF_X1 reg_mem_reg_94__6_ ( .D(n8996), .CK(clk), .Q(reg_mem[1294]) );
  DFF_X1 reg_mem_reg_94__5_ ( .D(n8995), .CK(clk), .Q(reg_mem[1293]) );
  DFF_X1 reg_mem_reg_94__4_ ( .D(n8994), .CK(clk), .Q(reg_mem[1292]) );
  DFF_X1 reg_mem_reg_94__3_ ( .D(n8993), .CK(clk), .Q(reg_mem[1291]) );
  DFF_X1 reg_mem_reg_94__2_ ( .D(n8992), .CK(clk), .Q(reg_mem[1290]) );
  DFF_X1 reg_mem_reg_94__1_ ( .D(n8991), .CK(clk), .Q(reg_mem[1289]) );
  DFF_X1 reg_mem_reg_94__0_ ( .D(n8990), .CK(clk), .Q(reg_mem[1288]) );
  DFF_X1 reg_mem_reg_95__7_ ( .D(n7268), .CK(clk), .Q(reg_mem[1287]) );
  DFF_X1 reg_mem_reg_95__6_ ( .D(n7267), .CK(clk), .Q(reg_mem[1286]) );
  DFF_X1 reg_mem_reg_95__5_ ( .D(n7266), .CK(clk), .Q(reg_mem[1285]) );
  DFF_X1 reg_mem_reg_95__4_ ( .D(n7265), .CK(clk), .Q(reg_mem[1284]) );
  DFF_X1 reg_mem_reg_95__3_ ( .D(n7264), .CK(clk), .Q(reg_mem[1283]) );
  DFF_X1 reg_mem_reg_95__2_ ( .D(n7263), .CK(clk), .Q(reg_mem[1282]) );
  DFF_X1 reg_mem_reg_95__1_ ( .D(n7262), .CK(clk), .Q(reg_mem[1281]) );
  DFF_X1 reg_mem_reg_95__0_ ( .D(n7261), .CK(clk), .Q(reg_mem[1280]) );
  DFF_X1 reg_mem_reg_96__7_ ( .D(n7998), .CK(clk), .Q(reg_mem[1279]) );
  DFF_X1 reg_mem_reg_96__6_ ( .D(n7997), .CK(clk), .Q(reg_mem[1278]) );
  DFF_X1 reg_mem_reg_96__5_ ( .D(n7996), .CK(clk), .Q(reg_mem[1277]) );
  DFF_X1 reg_mem_reg_96__4_ ( .D(n7995), .CK(clk), .Q(reg_mem[1276]) );
  DFF_X1 reg_mem_reg_96__3_ ( .D(n7994), .CK(clk), .Q(reg_mem[1275]) );
  DFF_X1 reg_mem_reg_96__2_ ( .D(n7993), .CK(clk), .Q(reg_mem[1274]) );
  DFF_X1 reg_mem_reg_96__1_ ( .D(n7992), .CK(clk), .Q(reg_mem[1273]) );
  DFF_X1 reg_mem_reg_96__0_ ( .D(n7991), .CK(clk), .Q(reg_mem[1272]) );
  DFF_X1 reg_mem_reg_97__7_ ( .D(n7421), .CK(clk), .Q(reg_mem[1271]) );
  DFF_X1 reg_mem_reg_97__6_ ( .D(n7420), .CK(clk), .Q(reg_mem[1270]) );
  DFF_X1 reg_mem_reg_97__5_ ( .D(n7419), .CK(clk), .Q(reg_mem[1269]) );
  DFF_X1 reg_mem_reg_97__4_ ( .D(n7418), .CK(clk), .Q(reg_mem[1268]) );
  DFF_X1 reg_mem_reg_97__3_ ( .D(n7417), .CK(clk), .Q(reg_mem[1267]) );
  DFF_X1 reg_mem_reg_97__2_ ( .D(n7416), .CK(clk), .Q(reg_mem[1266]) );
  DFF_X1 reg_mem_reg_97__1_ ( .D(n7415), .CK(clk), .Q(reg_mem[1265]) );
  DFF_X1 reg_mem_reg_97__0_ ( .D(n7414), .CK(clk), .Q(reg_mem[1264]) );
  DFF_X1 reg_mem_reg_98__7_ ( .D(n8574), .CK(clk), .Q(reg_mem[1263]) );
  DFF_X1 reg_mem_reg_98__6_ ( .D(n8573), .CK(clk), .Q(reg_mem[1262]) );
  DFF_X1 reg_mem_reg_98__5_ ( .D(n8572), .CK(clk), .Q(reg_mem[1261]) );
  DFF_X1 reg_mem_reg_98__4_ ( .D(n8571), .CK(clk), .Q(reg_mem[1260]) );
  DFF_X1 reg_mem_reg_98__3_ ( .D(n8570), .CK(clk), .Q(reg_mem[1259]) );
  DFF_X1 reg_mem_reg_98__2_ ( .D(n8569), .CK(clk), .Q(reg_mem[1258]) );
  DFF_X1 reg_mem_reg_98__1_ ( .D(n8568), .CK(clk), .Q(reg_mem[1257]) );
  DFF_X1 reg_mem_reg_98__0_ ( .D(n8567), .CK(clk), .Q(reg_mem[1256]) );
  DFF_X1 reg_mem_reg_99__7_ ( .D(n6845), .CK(clk), .Q(reg_mem[1255]) );
  DFF_X1 reg_mem_reg_99__6_ ( .D(n6844), .CK(clk), .Q(reg_mem[1254]) );
  DFF_X1 reg_mem_reg_99__5_ ( .D(n6843), .CK(clk), .Q(reg_mem[1253]) );
  DFF_X1 reg_mem_reg_99__4_ ( .D(n6842), .CK(clk), .Q(reg_mem[1252]) );
  DFF_X1 reg_mem_reg_99__3_ ( .D(n6841), .CK(clk), .Q(reg_mem[1251]) );
  DFF_X1 reg_mem_reg_99__2_ ( .D(n6840), .CK(clk), .Q(reg_mem[1250]) );
  DFF_X1 reg_mem_reg_99__1_ ( .D(n6839), .CK(clk), .Q(reg_mem[1249]) );
  DFF_X1 reg_mem_reg_99__0_ ( .D(n6838), .CK(clk), .Q(reg_mem[1248]) );
  DFF_X1 reg_mem_reg_100__7_ ( .D(n8142), .CK(clk), .Q(reg_mem[1247]) );
  DFF_X1 reg_mem_reg_100__6_ ( .D(n8141), .CK(clk), .Q(reg_mem[1246]) );
  DFF_X1 reg_mem_reg_100__5_ ( .D(n8140), .CK(clk), .Q(reg_mem[1245]) );
  DFF_X1 reg_mem_reg_100__4_ ( .D(n8139), .CK(clk), .Q(reg_mem[1244]) );
  DFF_X1 reg_mem_reg_100__3_ ( .D(n8138), .CK(clk), .Q(reg_mem[1243]) );
  DFF_X1 reg_mem_reg_100__2_ ( .D(n8137), .CK(clk), .Q(reg_mem[1242]) );
  DFF_X1 reg_mem_reg_100__1_ ( .D(n8136), .CK(clk), .Q(reg_mem[1241]) );
  DFF_X1 reg_mem_reg_100__0_ ( .D(n8135), .CK(clk), .Q(reg_mem[1240]) );
  DFF_X1 reg_mem_reg_101__7_ ( .D(n7565), .CK(clk), .Q(reg_mem[1239]) );
  DFF_X1 reg_mem_reg_101__6_ ( .D(n7564), .CK(clk), .Q(reg_mem[1238]) );
  DFF_X1 reg_mem_reg_101__5_ ( .D(n7563), .CK(clk), .Q(reg_mem[1237]) );
  DFF_X1 reg_mem_reg_101__4_ ( .D(n7562), .CK(clk), .Q(reg_mem[1236]) );
  DFF_X1 reg_mem_reg_101__3_ ( .D(n7561), .CK(clk), .Q(reg_mem[1235]) );
  DFF_X1 reg_mem_reg_101__2_ ( .D(n7560), .CK(clk), .Q(reg_mem[1234]) );
  DFF_X1 reg_mem_reg_101__1_ ( .D(n7559), .CK(clk), .Q(reg_mem[1233]) );
  DFF_X1 reg_mem_reg_101__0_ ( .D(n7558), .CK(clk), .Q(reg_mem[1232]) );
  DFF_X1 reg_mem_reg_102__7_ ( .D(n8718), .CK(clk), .Q(reg_mem[1231]) );
  DFF_X1 reg_mem_reg_102__6_ ( .D(n8717), .CK(clk), .Q(reg_mem[1230]) );
  DFF_X1 reg_mem_reg_102__5_ ( .D(n8716), .CK(clk), .Q(reg_mem[1229]) );
  DFF_X1 reg_mem_reg_102__4_ ( .D(n8715), .CK(clk), .Q(reg_mem[1228]) );
  DFF_X1 reg_mem_reg_102__3_ ( .D(n8714), .CK(clk), .Q(reg_mem[1227]) );
  DFF_X1 reg_mem_reg_102__2_ ( .D(n8713), .CK(clk), .Q(reg_mem[1226]) );
  DFF_X1 reg_mem_reg_102__1_ ( .D(n8712), .CK(clk), .Q(reg_mem[1225]) );
  DFF_X1 reg_mem_reg_102__0_ ( .D(n8711), .CK(clk), .Q(reg_mem[1224]) );
  DFF_X1 reg_mem_reg_103__7_ ( .D(n6989), .CK(clk), .Q(reg_mem[1223]) );
  DFF_X1 reg_mem_reg_103__6_ ( .D(n6988), .CK(clk), .Q(reg_mem[1222]) );
  DFF_X1 reg_mem_reg_103__5_ ( .D(n6987), .CK(clk), .Q(reg_mem[1221]) );
  DFF_X1 reg_mem_reg_103__4_ ( .D(n6986), .CK(clk), .Q(reg_mem[1220]) );
  DFF_X1 reg_mem_reg_103__3_ ( .D(n6985), .CK(clk), .Q(reg_mem[1219]) );
  DFF_X1 reg_mem_reg_103__2_ ( .D(n6984), .CK(clk), .Q(reg_mem[1218]) );
  DFF_X1 reg_mem_reg_103__1_ ( .D(n6983), .CK(clk), .Q(reg_mem[1217]) );
  DFF_X1 reg_mem_reg_103__0_ ( .D(n6982), .CK(clk), .Q(reg_mem[1216]) );
  DFF_X1 reg_mem_reg_104__7_ ( .D(n8286), .CK(clk), .Q(reg_mem[1215]) );
  DFF_X1 reg_mem_reg_104__6_ ( .D(n8285), .CK(clk), .Q(reg_mem[1214]) );
  DFF_X1 reg_mem_reg_104__5_ ( .D(n8284), .CK(clk), .Q(reg_mem[1213]) );
  DFF_X1 reg_mem_reg_104__4_ ( .D(n8283), .CK(clk), .Q(reg_mem[1212]) );
  DFF_X1 reg_mem_reg_104__3_ ( .D(n8282), .CK(clk), .Q(reg_mem[1211]) );
  DFF_X1 reg_mem_reg_104__2_ ( .D(n8281), .CK(clk), .Q(reg_mem[1210]) );
  DFF_X1 reg_mem_reg_104__1_ ( .D(n8280), .CK(clk), .Q(reg_mem[1209]) );
  DFF_X1 reg_mem_reg_104__0_ ( .D(n8279), .CK(clk), .Q(reg_mem[1208]) );
  DFF_X1 reg_mem_reg_105__7_ ( .D(n7709), .CK(clk), .Q(reg_mem[1207]) );
  DFF_X1 reg_mem_reg_105__6_ ( .D(n7708), .CK(clk), .Q(reg_mem[1206]) );
  DFF_X1 reg_mem_reg_105__5_ ( .D(n7707), .CK(clk), .Q(reg_mem[1205]) );
  DFF_X1 reg_mem_reg_105__4_ ( .D(n7706), .CK(clk), .Q(reg_mem[1204]) );
  DFF_X1 reg_mem_reg_105__3_ ( .D(n7705), .CK(clk), .Q(reg_mem[1203]) );
  DFF_X1 reg_mem_reg_105__2_ ( .D(n7704), .CK(clk), .Q(reg_mem[1202]) );
  DFF_X1 reg_mem_reg_105__1_ ( .D(n7703), .CK(clk), .Q(reg_mem[1201]) );
  DFF_X1 reg_mem_reg_105__0_ ( .D(n7702), .CK(clk), .Q(reg_mem[1200]) );
  DFF_X1 reg_mem_reg_106__7_ ( .D(n8862), .CK(clk), .Q(reg_mem[1199]) );
  DFF_X1 reg_mem_reg_106__6_ ( .D(n8861), .CK(clk), .Q(reg_mem[1198]) );
  DFF_X1 reg_mem_reg_106__5_ ( .D(n8860), .CK(clk), .Q(reg_mem[1197]) );
  DFF_X1 reg_mem_reg_106__4_ ( .D(n8859), .CK(clk), .Q(reg_mem[1196]) );
  DFF_X1 reg_mem_reg_106__3_ ( .D(n8858), .CK(clk), .Q(reg_mem[1195]) );
  DFF_X1 reg_mem_reg_106__2_ ( .D(n8857), .CK(clk), .Q(reg_mem[1194]) );
  DFF_X1 reg_mem_reg_106__1_ ( .D(n8856), .CK(clk), .Q(reg_mem[1193]) );
  DFF_X1 reg_mem_reg_106__0_ ( .D(n8855), .CK(clk), .Q(reg_mem[1192]) );
  DFF_X1 reg_mem_reg_107__7_ ( .D(n7133), .CK(clk), .Q(reg_mem[1191]) );
  DFF_X1 reg_mem_reg_107__6_ ( .D(n7132), .CK(clk), .Q(reg_mem[1190]) );
  DFF_X1 reg_mem_reg_107__5_ ( .D(n7131), .CK(clk), .Q(reg_mem[1189]) );
  DFF_X1 reg_mem_reg_107__4_ ( .D(n7130), .CK(clk), .Q(reg_mem[1188]) );
  DFF_X1 reg_mem_reg_107__3_ ( .D(n7129), .CK(clk), .Q(reg_mem[1187]) );
  DFF_X1 reg_mem_reg_107__2_ ( .D(n7128), .CK(clk), .Q(reg_mem[1186]) );
  DFF_X1 reg_mem_reg_107__1_ ( .D(n7127), .CK(clk), .Q(reg_mem[1185]) );
  DFF_X1 reg_mem_reg_107__0_ ( .D(n7126), .CK(clk), .Q(reg_mem[1184]) );
  DFF_X1 reg_mem_reg_108__7_ ( .D(n8430), .CK(clk), .Q(reg_mem[1183]) );
  DFF_X1 reg_mem_reg_108__6_ ( .D(n8429), .CK(clk), .Q(reg_mem[1182]) );
  DFF_X1 reg_mem_reg_108__5_ ( .D(n8428), .CK(clk), .Q(reg_mem[1181]) );
  DFF_X1 reg_mem_reg_108__4_ ( .D(n8427), .CK(clk), .Q(reg_mem[1180]) );
  DFF_X1 reg_mem_reg_108__3_ ( .D(n8426), .CK(clk), .Q(reg_mem[1179]) );
  DFF_X1 reg_mem_reg_108__2_ ( .D(n8425), .CK(clk), .Q(reg_mem[1178]) );
  DFF_X1 reg_mem_reg_108__1_ ( .D(n8424), .CK(clk), .Q(reg_mem[1177]) );
  DFF_X1 reg_mem_reg_108__0_ ( .D(n8423), .CK(clk), .Q(reg_mem[1176]) );
  DFF_X1 reg_mem_reg_109__7_ ( .D(n7853), .CK(clk), .Q(reg_mem[1175]) );
  DFF_X1 reg_mem_reg_109__6_ ( .D(n7852), .CK(clk), .Q(reg_mem[1174]) );
  DFF_X1 reg_mem_reg_109__5_ ( .D(n7851), .CK(clk), .Q(reg_mem[1173]) );
  DFF_X1 reg_mem_reg_109__4_ ( .D(n7850), .CK(clk), .Q(reg_mem[1172]) );
  DFF_X1 reg_mem_reg_109__3_ ( .D(n7849), .CK(clk), .Q(reg_mem[1171]) );
  DFF_X1 reg_mem_reg_109__2_ ( .D(n7848), .CK(clk), .Q(reg_mem[1170]) );
  DFF_X1 reg_mem_reg_109__1_ ( .D(n7847), .CK(clk), .Q(reg_mem[1169]) );
  DFF_X1 reg_mem_reg_109__0_ ( .D(n7846), .CK(clk), .Q(reg_mem[1168]) );
  DFF_X1 reg_mem_reg_110__7_ ( .D(n9006), .CK(clk), .Q(reg_mem[1167]) );
  DFF_X1 reg_mem_reg_110__6_ ( .D(n9005), .CK(clk), .Q(reg_mem[1166]) );
  DFF_X1 reg_mem_reg_110__5_ ( .D(n9004), .CK(clk), .Q(reg_mem[1165]) );
  DFF_X1 reg_mem_reg_110__4_ ( .D(n9003), .CK(clk), .Q(reg_mem[1164]) );
  DFF_X1 reg_mem_reg_110__3_ ( .D(n9002), .CK(clk), .Q(reg_mem[1163]) );
  DFF_X1 reg_mem_reg_110__2_ ( .D(n9001), .CK(clk), .Q(reg_mem[1162]) );
  DFF_X1 reg_mem_reg_110__1_ ( .D(n9000), .CK(clk), .Q(reg_mem[1161]) );
  DFF_X1 reg_mem_reg_110__0_ ( .D(n8999), .CK(clk), .Q(reg_mem[1160]) );
  DFF_X1 reg_mem_reg_111__7_ ( .D(n7277), .CK(clk), .Q(reg_mem[1159]) );
  DFF_X1 reg_mem_reg_111__6_ ( .D(n7276), .CK(clk), .Q(reg_mem[1158]) );
  DFF_X1 reg_mem_reg_111__5_ ( .D(n7275), .CK(clk), .Q(reg_mem[1157]) );
  DFF_X1 reg_mem_reg_111__4_ ( .D(n7274), .CK(clk), .Q(reg_mem[1156]) );
  DFF_X1 reg_mem_reg_111__3_ ( .D(n7273), .CK(clk), .Q(reg_mem[1155]) );
  DFF_X1 reg_mem_reg_111__2_ ( .D(n7272), .CK(clk), .Q(reg_mem[1154]) );
  DFF_X1 reg_mem_reg_111__1_ ( .D(n7271), .CK(clk), .Q(reg_mem[1153]) );
  DFF_X1 reg_mem_reg_111__0_ ( .D(n7270), .CK(clk), .Q(reg_mem[1152]) );
  DFF_X1 reg_mem_reg_112__7_ ( .D(n8007), .CK(clk), .Q(reg_mem[1151]) );
  DFF_X1 reg_mem_reg_112__6_ ( .D(n8006), .CK(clk), .Q(reg_mem[1150]) );
  DFF_X1 reg_mem_reg_112__5_ ( .D(n8005), .CK(clk), .Q(reg_mem[1149]) );
  DFF_X1 reg_mem_reg_112__4_ ( .D(n8004), .CK(clk), .Q(reg_mem[1148]) );
  DFF_X1 reg_mem_reg_112__3_ ( .D(n8003), .CK(clk), .Q(reg_mem[1147]) );
  DFF_X1 reg_mem_reg_112__2_ ( .D(n8002), .CK(clk), .Q(reg_mem[1146]) );
  DFF_X1 reg_mem_reg_112__1_ ( .D(n8001), .CK(clk), .Q(reg_mem[1145]) );
  DFF_X1 reg_mem_reg_112__0_ ( .D(n8000), .CK(clk), .Q(reg_mem[1144]) );
  DFF_X1 reg_mem_reg_113__7_ ( .D(n7430), .CK(clk), .Q(reg_mem[1143]) );
  DFF_X1 reg_mem_reg_113__6_ ( .D(n7429), .CK(clk), .Q(reg_mem[1142]) );
  DFF_X1 reg_mem_reg_113__5_ ( .D(n7428), .CK(clk), .Q(reg_mem[1141]) );
  DFF_X1 reg_mem_reg_113__4_ ( .D(n7427), .CK(clk), .Q(reg_mem[1140]) );
  DFF_X1 reg_mem_reg_113__3_ ( .D(n7426), .CK(clk), .Q(reg_mem[1139]) );
  DFF_X1 reg_mem_reg_113__2_ ( .D(n7425), .CK(clk), .Q(reg_mem[1138]) );
  DFF_X1 reg_mem_reg_113__1_ ( .D(n7424), .CK(clk), .Q(reg_mem[1137]) );
  DFF_X1 reg_mem_reg_113__0_ ( .D(n7423), .CK(clk), .Q(reg_mem[1136]) );
  DFF_X1 reg_mem_reg_114__7_ ( .D(n8583), .CK(clk), .Q(reg_mem[1135]) );
  DFF_X1 reg_mem_reg_114__6_ ( .D(n8582), .CK(clk), .Q(reg_mem[1134]) );
  DFF_X1 reg_mem_reg_114__5_ ( .D(n8581), .CK(clk), .Q(reg_mem[1133]) );
  DFF_X1 reg_mem_reg_114__4_ ( .D(n8580), .CK(clk), .Q(reg_mem[1132]) );
  DFF_X1 reg_mem_reg_114__3_ ( .D(n8579), .CK(clk), .Q(reg_mem[1131]) );
  DFF_X1 reg_mem_reg_114__2_ ( .D(n8578), .CK(clk), .Q(reg_mem[1130]) );
  DFF_X1 reg_mem_reg_114__1_ ( .D(n8577), .CK(clk), .Q(reg_mem[1129]) );
  DFF_X1 reg_mem_reg_114__0_ ( .D(n8576), .CK(clk), .Q(reg_mem[1128]) );
  DFF_X1 reg_mem_reg_115__7_ ( .D(n6854), .CK(clk), .Q(reg_mem[1127]) );
  DFF_X1 reg_mem_reg_115__6_ ( .D(n6853), .CK(clk), .Q(reg_mem[1126]) );
  DFF_X1 reg_mem_reg_115__5_ ( .D(n6852), .CK(clk), .Q(reg_mem[1125]) );
  DFF_X1 reg_mem_reg_115__4_ ( .D(n6851), .CK(clk), .Q(reg_mem[1124]) );
  DFF_X1 reg_mem_reg_115__3_ ( .D(n6850), .CK(clk), .Q(reg_mem[1123]) );
  DFF_X1 reg_mem_reg_115__2_ ( .D(n6849), .CK(clk), .Q(reg_mem[1122]) );
  DFF_X1 reg_mem_reg_115__1_ ( .D(n6848), .CK(clk), .Q(reg_mem[1121]) );
  DFF_X1 reg_mem_reg_115__0_ ( .D(n6847), .CK(clk), .Q(reg_mem[1120]) );
  DFF_X1 reg_mem_reg_116__7_ ( .D(n8151), .CK(clk), .Q(reg_mem[1119]) );
  DFF_X1 reg_mem_reg_116__6_ ( .D(n8150), .CK(clk), .Q(reg_mem[1118]) );
  DFF_X1 reg_mem_reg_116__5_ ( .D(n8149), .CK(clk), .Q(reg_mem[1117]) );
  DFF_X1 reg_mem_reg_116__4_ ( .D(n8148), .CK(clk), .Q(reg_mem[1116]) );
  DFF_X1 reg_mem_reg_116__3_ ( .D(n8147), .CK(clk), .Q(reg_mem[1115]) );
  DFF_X1 reg_mem_reg_116__2_ ( .D(n8146), .CK(clk), .Q(reg_mem[1114]) );
  DFF_X1 reg_mem_reg_116__1_ ( .D(n8145), .CK(clk), .Q(reg_mem[1113]) );
  DFF_X1 reg_mem_reg_116__0_ ( .D(n8144), .CK(clk), .Q(reg_mem[1112]) );
  DFF_X1 reg_mem_reg_117__7_ ( .D(n7574), .CK(clk), .Q(reg_mem[1111]) );
  DFF_X1 reg_mem_reg_117__6_ ( .D(n7573), .CK(clk), .Q(reg_mem[1110]) );
  DFF_X1 reg_mem_reg_117__5_ ( .D(n7572), .CK(clk), .Q(reg_mem[1109]) );
  DFF_X1 reg_mem_reg_117__4_ ( .D(n7571), .CK(clk), .Q(reg_mem[1108]) );
  DFF_X1 reg_mem_reg_117__3_ ( .D(n7570), .CK(clk), .Q(reg_mem[1107]) );
  DFF_X1 reg_mem_reg_117__2_ ( .D(n7569), .CK(clk), .Q(reg_mem[1106]) );
  DFF_X1 reg_mem_reg_117__1_ ( .D(n7568), .CK(clk), .Q(reg_mem[1105]) );
  DFF_X1 reg_mem_reg_117__0_ ( .D(n7567), .CK(clk), .Q(reg_mem[1104]) );
  DFF_X1 reg_mem_reg_118__7_ ( .D(n8727), .CK(clk), .Q(reg_mem[1103]) );
  DFF_X1 reg_mem_reg_118__6_ ( .D(n8726), .CK(clk), .Q(reg_mem[1102]) );
  DFF_X1 reg_mem_reg_118__5_ ( .D(n8725), .CK(clk), .Q(reg_mem[1101]) );
  DFF_X1 reg_mem_reg_118__4_ ( .D(n8724), .CK(clk), .Q(reg_mem[1100]) );
  DFF_X1 reg_mem_reg_118__3_ ( .D(n8723), .CK(clk), .Q(reg_mem[1099]) );
  DFF_X1 reg_mem_reg_118__2_ ( .D(n8722), .CK(clk), .Q(reg_mem[1098]) );
  DFF_X1 reg_mem_reg_118__1_ ( .D(n8721), .CK(clk), .Q(reg_mem[1097]) );
  DFF_X1 reg_mem_reg_118__0_ ( .D(n8720), .CK(clk), .Q(reg_mem[1096]) );
  DFF_X1 reg_mem_reg_119__7_ ( .D(n6998), .CK(clk), .Q(reg_mem[1095]) );
  DFF_X1 reg_mem_reg_119__6_ ( .D(n6997), .CK(clk), .Q(reg_mem[1094]) );
  DFF_X1 reg_mem_reg_119__5_ ( .D(n6996), .CK(clk), .Q(reg_mem[1093]) );
  DFF_X1 reg_mem_reg_119__4_ ( .D(n6995), .CK(clk), .Q(reg_mem[1092]) );
  DFF_X1 reg_mem_reg_119__3_ ( .D(n6994), .CK(clk), .Q(reg_mem[1091]) );
  DFF_X1 reg_mem_reg_119__2_ ( .D(n6993), .CK(clk), .Q(reg_mem[1090]) );
  DFF_X1 reg_mem_reg_119__1_ ( .D(n6992), .CK(clk), .Q(reg_mem[1089]) );
  DFF_X1 reg_mem_reg_119__0_ ( .D(n6991), .CK(clk), .Q(reg_mem[1088]) );
  DFF_X1 reg_mem_reg_120__7_ ( .D(n8295), .CK(clk), .Q(reg_mem[1087]) );
  DFF_X1 reg_mem_reg_120__6_ ( .D(n8294), .CK(clk), .Q(reg_mem[1086]) );
  DFF_X1 reg_mem_reg_120__5_ ( .D(n8293), .CK(clk), .Q(reg_mem[1085]) );
  DFF_X1 reg_mem_reg_120__4_ ( .D(n8292), .CK(clk), .Q(reg_mem[1084]) );
  DFF_X1 reg_mem_reg_120__3_ ( .D(n8291), .CK(clk), .Q(reg_mem[1083]) );
  DFF_X1 reg_mem_reg_120__2_ ( .D(n8290), .CK(clk), .Q(reg_mem[1082]) );
  DFF_X1 reg_mem_reg_120__1_ ( .D(n8289), .CK(clk), .Q(reg_mem[1081]) );
  DFF_X1 reg_mem_reg_120__0_ ( .D(n8288), .CK(clk), .Q(reg_mem[1080]) );
  DFF_X1 reg_mem_reg_121__7_ ( .D(n7718), .CK(clk), .Q(reg_mem[1079]) );
  DFF_X1 reg_mem_reg_121__6_ ( .D(n7717), .CK(clk), .Q(reg_mem[1078]) );
  DFF_X1 reg_mem_reg_121__5_ ( .D(n7716), .CK(clk), .Q(reg_mem[1077]) );
  DFF_X1 reg_mem_reg_121__4_ ( .D(n7715), .CK(clk), .Q(reg_mem[1076]) );
  DFF_X1 reg_mem_reg_121__3_ ( .D(n7714), .CK(clk), .Q(reg_mem[1075]) );
  DFF_X1 reg_mem_reg_121__2_ ( .D(n7713), .CK(clk), .Q(reg_mem[1074]) );
  DFF_X1 reg_mem_reg_121__1_ ( .D(n7712), .CK(clk), .Q(reg_mem[1073]) );
  DFF_X1 reg_mem_reg_121__0_ ( .D(n7711), .CK(clk), .Q(reg_mem[1072]) );
  DFF_X1 reg_mem_reg_122__7_ ( .D(n8871), .CK(clk), .Q(reg_mem[1071]) );
  DFF_X1 reg_mem_reg_122__6_ ( .D(n8870), .CK(clk), .Q(reg_mem[1070]) );
  DFF_X1 reg_mem_reg_122__5_ ( .D(n8869), .CK(clk), .Q(reg_mem[1069]) );
  DFF_X1 reg_mem_reg_122__4_ ( .D(n8868), .CK(clk), .Q(reg_mem[1068]) );
  DFF_X1 reg_mem_reg_122__3_ ( .D(n8867), .CK(clk), .Q(reg_mem[1067]) );
  DFF_X1 reg_mem_reg_122__2_ ( .D(n8866), .CK(clk), .Q(reg_mem[1066]) );
  DFF_X1 reg_mem_reg_122__1_ ( .D(n8865), .CK(clk), .Q(reg_mem[1065]) );
  DFF_X1 reg_mem_reg_122__0_ ( .D(n8864), .CK(clk), .Q(reg_mem[1064]) );
  DFF_X1 reg_mem_reg_123__7_ ( .D(n7142), .CK(clk), .Q(reg_mem[1063]) );
  DFF_X1 reg_mem_reg_123__6_ ( .D(n7141), .CK(clk), .Q(reg_mem[1062]) );
  DFF_X1 reg_mem_reg_123__5_ ( .D(n7140), .CK(clk), .Q(reg_mem[1061]) );
  DFF_X1 reg_mem_reg_123__4_ ( .D(n7139), .CK(clk), .Q(reg_mem[1060]) );
  DFF_X1 reg_mem_reg_123__3_ ( .D(n7138), .CK(clk), .Q(reg_mem[1059]) );
  DFF_X1 reg_mem_reg_123__2_ ( .D(n7137), .CK(clk), .Q(reg_mem[1058]) );
  DFF_X1 reg_mem_reg_123__1_ ( .D(n7136), .CK(clk), .Q(reg_mem[1057]) );
  DFF_X1 reg_mem_reg_123__0_ ( .D(n7135), .CK(clk), .Q(reg_mem[1056]) );
  DFF_X1 reg_mem_reg_124__7_ ( .D(n8439), .CK(clk), .Q(reg_mem[1055]) );
  DFF_X1 reg_mem_reg_124__6_ ( .D(n8438), .CK(clk), .Q(reg_mem[1054]) );
  DFF_X1 reg_mem_reg_124__5_ ( .D(n8437), .CK(clk), .Q(reg_mem[1053]) );
  DFF_X1 reg_mem_reg_124__4_ ( .D(n8436), .CK(clk), .Q(reg_mem[1052]) );
  DFF_X1 reg_mem_reg_124__3_ ( .D(n8435), .CK(clk), .Q(reg_mem[1051]) );
  DFF_X1 reg_mem_reg_124__2_ ( .D(n8434), .CK(clk), .Q(reg_mem[1050]) );
  DFF_X1 reg_mem_reg_124__1_ ( .D(n8433), .CK(clk), .Q(reg_mem[1049]) );
  DFF_X1 reg_mem_reg_124__0_ ( .D(n8432), .CK(clk), .Q(reg_mem[1048]) );
  DFF_X1 reg_mem_reg_125__7_ ( .D(n7862), .CK(clk), .Q(reg_mem[1047]) );
  DFF_X1 reg_mem_reg_125__6_ ( .D(n7861), .CK(clk), .Q(reg_mem[1046]) );
  DFF_X1 reg_mem_reg_125__5_ ( .D(n7860), .CK(clk), .Q(reg_mem[1045]) );
  DFF_X1 reg_mem_reg_125__4_ ( .D(n7859), .CK(clk), .Q(reg_mem[1044]) );
  DFF_X1 reg_mem_reg_125__3_ ( .D(n7858), .CK(clk), .Q(reg_mem[1043]) );
  DFF_X1 reg_mem_reg_125__2_ ( .D(n7857), .CK(clk), .Q(reg_mem[1042]) );
  DFF_X1 reg_mem_reg_125__1_ ( .D(n7856), .CK(clk), .Q(reg_mem[1041]) );
  DFF_X1 reg_mem_reg_125__0_ ( .D(n7855), .CK(clk), .Q(reg_mem[1040]) );
  DFF_X1 reg_mem_reg_126__7_ ( .D(n9015), .CK(clk), .Q(reg_mem[1039]) );
  DFF_X1 reg_mem_reg_126__6_ ( .D(n9014), .CK(clk), .Q(reg_mem[1038]) );
  DFF_X1 reg_mem_reg_126__5_ ( .D(n9013), .CK(clk), .Q(reg_mem[1037]) );
  DFF_X1 reg_mem_reg_126__4_ ( .D(n9012), .CK(clk), .Q(reg_mem[1036]) );
  DFF_X1 reg_mem_reg_126__3_ ( .D(n9011), .CK(clk), .Q(reg_mem[1035]) );
  DFF_X1 reg_mem_reg_126__2_ ( .D(n9010), .CK(clk), .Q(reg_mem[1034]) );
  DFF_X1 reg_mem_reg_126__1_ ( .D(n9009), .CK(clk), .Q(reg_mem[1033]) );
  DFF_X1 reg_mem_reg_126__0_ ( .D(n9008), .CK(clk), .Q(reg_mem[1032]) );
  DFF_X1 reg_mem_reg_127__7_ ( .D(n7286), .CK(clk), .Q(reg_mem[1031]) );
  DFF_X1 reg_mem_reg_127__6_ ( .D(n7285), .CK(clk), .Q(reg_mem[1030]) );
  DFF_X1 reg_mem_reg_127__5_ ( .D(n7284), .CK(clk), .Q(reg_mem[1029]) );
  DFF_X1 reg_mem_reg_127__4_ ( .D(n7283), .CK(clk), .Q(reg_mem[1028]) );
  DFF_X1 reg_mem_reg_127__3_ ( .D(n7282), .CK(clk), .Q(reg_mem[1027]) );
  DFF_X1 reg_mem_reg_127__2_ ( .D(n7281), .CK(clk), .Q(reg_mem[1026]) );
  DFF_X1 reg_mem_reg_127__1_ ( .D(n7280), .CK(clk), .Q(reg_mem[1025]) );
  DFF_X1 reg_mem_reg_127__0_ ( .D(n7279), .CK(clk), .Q(reg_mem[1024]) );
  DFF_X1 reg_mem_reg_128__7_ ( .D(n8016), .CK(clk), .Q(reg_mem[1023]) );
  DFF_X1 reg_mem_reg_128__6_ ( .D(n8015), .CK(clk), .Q(reg_mem[1022]) );
  DFF_X1 reg_mem_reg_128__5_ ( .D(n8014), .CK(clk), .Q(reg_mem[1021]) );
  DFF_X1 reg_mem_reg_128__4_ ( .D(n8013), .CK(clk), .Q(reg_mem[1020]) );
  DFF_X1 reg_mem_reg_128__3_ ( .D(n8012), .CK(clk), .Q(reg_mem[1019]) );
  DFF_X1 reg_mem_reg_128__2_ ( .D(n8011), .CK(clk), .Q(reg_mem[1018]) );
  DFF_X1 reg_mem_reg_128__1_ ( .D(n8010), .CK(clk), .Q(reg_mem[1017]) );
  DFF_X1 reg_mem_reg_128__0_ ( .D(n8009), .CK(clk), .Q(reg_mem[1016]) );
  DFF_X1 reg_mem_reg_129__7_ ( .D(n7439), .CK(clk), .Q(reg_mem[1015]) );
  DFF_X1 reg_mem_reg_129__6_ ( .D(n7438), .CK(clk), .Q(reg_mem[1014]) );
  DFF_X1 reg_mem_reg_129__5_ ( .D(n7437), .CK(clk), .Q(reg_mem[1013]) );
  DFF_X1 reg_mem_reg_129__4_ ( .D(n7436), .CK(clk), .Q(reg_mem[1012]) );
  DFF_X1 reg_mem_reg_129__3_ ( .D(n7435), .CK(clk), .Q(reg_mem[1011]) );
  DFF_X1 reg_mem_reg_129__2_ ( .D(n7434), .CK(clk), .Q(reg_mem[1010]) );
  DFF_X1 reg_mem_reg_129__1_ ( .D(n7433), .CK(clk), .Q(reg_mem[1009]) );
  DFF_X1 reg_mem_reg_129__0_ ( .D(n7432), .CK(clk), .Q(reg_mem[1008]) );
  DFF_X1 reg_mem_reg_130__7_ ( .D(n8592), .CK(clk), .Q(reg_mem[1007]) );
  DFF_X1 reg_mem_reg_130__6_ ( .D(n8591), .CK(clk), .Q(reg_mem[1006]) );
  DFF_X1 reg_mem_reg_130__5_ ( .D(n8590), .CK(clk), .Q(reg_mem[1005]) );
  DFF_X1 reg_mem_reg_130__4_ ( .D(n8589), .CK(clk), .Q(reg_mem[1004]) );
  DFF_X1 reg_mem_reg_130__3_ ( .D(n8588), .CK(clk), .Q(reg_mem[1003]) );
  DFF_X1 reg_mem_reg_130__2_ ( .D(n8587), .CK(clk), .Q(reg_mem[1002]) );
  DFF_X1 reg_mem_reg_130__1_ ( .D(n8586), .CK(clk), .Q(reg_mem[1001]) );
  DFF_X1 reg_mem_reg_130__0_ ( .D(n8585), .CK(clk), .Q(reg_mem[1000]) );
  DFF_X1 reg_mem_reg_131__7_ ( .D(n6863), .CK(clk), .Q(reg_mem[999]) );
  DFF_X1 reg_mem_reg_131__6_ ( .D(n6862), .CK(clk), .Q(reg_mem[998]) );
  DFF_X1 reg_mem_reg_131__5_ ( .D(n6861), .CK(clk), .Q(reg_mem[997]) );
  DFF_X1 reg_mem_reg_131__4_ ( .D(n6860), .CK(clk), .Q(reg_mem[996]) );
  DFF_X1 reg_mem_reg_131__3_ ( .D(n6859), .CK(clk), .Q(reg_mem[995]) );
  DFF_X1 reg_mem_reg_131__2_ ( .D(n6858), .CK(clk), .Q(reg_mem[994]) );
  DFF_X1 reg_mem_reg_131__1_ ( .D(n6857), .CK(clk), .Q(reg_mem[993]) );
  DFF_X1 reg_mem_reg_131__0_ ( .D(n6856), .CK(clk), .Q(reg_mem[992]) );
  DFF_X1 reg_mem_reg_132__7_ ( .D(n8160), .CK(clk), .Q(reg_mem[991]) );
  DFF_X1 reg_mem_reg_132__6_ ( .D(n8159), .CK(clk), .Q(reg_mem[990]) );
  DFF_X1 reg_mem_reg_132__5_ ( .D(n8158), .CK(clk), .Q(reg_mem[989]) );
  DFF_X1 reg_mem_reg_132__4_ ( .D(n8157), .CK(clk), .Q(reg_mem[988]) );
  DFF_X1 reg_mem_reg_132__3_ ( .D(n8156), .CK(clk), .Q(reg_mem[987]) );
  DFF_X1 reg_mem_reg_132__2_ ( .D(n8155), .CK(clk), .Q(reg_mem[986]) );
  DFF_X1 reg_mem_reg_132__1_ ( .D(n8154), .CK(clk), .Q(reg_mem[985]) );
  DFF_X1 reg_mem_reg_132__0_ ( .D(n8153), .CK(clk), .Q(reg_mem[984]) );
  DFF_X1 reg_mem_reg_133__7_ ( .D(n7583), .CK(clk), .Q(reg_mem[983]) );
  DFF_X1 reg_mem_reg_133__6_ ( .D(n7582), .CK(clk), .Q(reg_mem[982]) );
  DFF_X1 reg_mem_reg_133__5_ ( .D(n7581), .CK(clk), .Q(reg_mem[981]) );
  DFF_X1 reg_mem_reg_133__4_ ( .D(n7580), .CK(clk), .Q(reg_mem[980]) );
  DFF_X1 reg_mem_reg_133__3_ ( .D(n7579), .CK(clk), .Q(reg_mem[979]) );
  DFF_X1 reg_mem_reg_133__2_ ( .D(n7578), .CK(clk), .Q(reg_mem[978]) );
  DFF_X1 reg_mem_reg_133__1_ ( .D(n7577), .CK(clk), .Q(reg_mem[977]) );
  DFF_X1 reg_mem_reg_133__0_ ( .D(n7576), .CK(clk), .Q(reg_mem[976]) );
  DFF_X1 reg_mem_reg_134__7_ ( .D(n8736), .CK(clk), .Q(reg_mem[975]) );
  DFF_X1 reg_mem_reg_134__6_ ( .D(n8735), .CK(clk), .Q(reg_mem[974]) );
  DFF_X1 reg_mem_reg_134__5_ ( .D(n8734), .CK(clk), .Q(reg_mem[973]) );
  DFF_X1 reg_mem_reg_134__4_ ( .D(n8733), .CK(clk), .Q(reg_mem[972]) );
  DFF_X1 reg_mem_reg_134__3_ ( .D(n8732), .CK(clk), .Q(reg_mem[971]) );
  DFF_X1 reg_mem_reg_134__2_ ( .D(n8731), .CK(clk), .Q(reg_mem[970]) );
  DFF_X1 reg_mem_reg_134__1_ ( .D(n8730), .CK(clk), .Q(reg_mem[969]) );
  DFF_X1 reg_mem_reg_134__0_ ( .D(n8729), .CK(clk), .Q(reg_mem[968]) );
  DFF_X1 reg_mem_reg_135__7_ ( .D(n7007), .CK(clk), .Q(reg_mem[967]) );
  DFF_X1 reg_mem_reg_135__6_ ( .D(n7006), .CK(clk), .Q(reg_mem[966]) );
  DFF_X1 reg_mem_reg_135__5_ ( .D(n7005), .CK(clk), .Q(reg_mem[965]) );
  DFF_X1 reg_mem_reg_135__4_ ( .D(n7004), .CK(clk), .Q(reg_mem[964]) );
  DFF_X1 reg_mem_reg_135__3_ ( .D(n7003), .CK(clk), .Q(reg_mem[963]) );
  DFF_X1 reg_mem_reg_135__2_ ( .D(n7002), .CK(clk), .Q(reg_mem[962]) );
  DFF_X1 reg_mem_reg_135__1_ ( .D(n7001), .CK(clk), .Q(reg_mem[961]) );
  DFF_X1 reg_mem_reg_135__0_ ( .D(n7000), .CK(clk), .Q(reg_mem[960]) );
  DFF_X1 reg_mem_reg_136__7_ ( .D(n8304), .CK(clk), .Q(reg_mem[959]) );
  DFF_X1 reg_mem_reg_136__6_ ( .D(n8303), .CK(clk), .Q(reg_mem[958]) );
  DFF_X1 reg_mem_reg_136__5_ ( .D(n8302), .CK(clk), .Q(reg_mem[957]) );
  DFF_X1 reg_mem_reg_136__4_ ( .D(n8301), .CK(clk), .Q(reg_mem[956]) );
  DFF_X1 reg_mem_reg_136__3_ ( .D(n8300), .CK(clk), .Q(reg_mem[955]) );
  DFF_X1 reg_mem_reg_136__2_ ( .D(n8299), .CK(clk), .Q(reg_mem[954]) );
  DFF_X1 reg_mem_reg_136__1_ ( .D(n8298), .CK(clk), .Q(reg_mem[953]) );
  DFF_X1 reg_mem_reg_136__0_ ( .D(n8297), .CK(clk), .Q(reg_mem[952]) );
  DFF_X1 reg_mem_reg_137__7_ ( .D(n7727), .CK(clk), .Q(reg_mem[951]) );
  DFF_X1 reg_mem_reg_137__6_ ( .D(n7726), .CK(clk), .Q(reg_mem[950]) );
  DFF_X1 reg_mem_reg_137__5_ ( .D(n7725), .CK(clk), .Q(reg_mem[949]) );
  DFF_X1 reg_mem_reg_137__4_ ( .D(n7724), .CK(clk), .Q(reg_mem[948]) );
  DFF_X1 reg_mem_reg_137__3_ ( .D(n7723), .CK(clk), .Q(reg_mem[947]) );
  DFF_X1 reg_mem_reg_137__2_ ( .D(n7722), .CK(clk), .Q(reg_mem[946]) );
  DFF_X1 reg_mem_reg_137__1_ ( .D(n7721), .CK(clk), .Q(reg_mem[945]) );
  DFF_X1 reg_mem_reg_137__0_ ( .D(n7720), .CK(clk), .Q(reg_mem[944]) );
  DFF_X1 reg_mem_reg_138__7_ ( .D(n8880), .CK(clk), .Q(reg_mem[943]) );
  DFF_X1 reg_mem_reg_138__6_ ( .D(n8879), .CK(clk), .Q(reg_mem[942]) );
  DFF_X1 reg_mem_reg_138__5_ ( .D(n8878), .CK(clk), .Q(reg_mem[941]) );
  DFF_X1 reg_mem_reg_138__4_ ( .D(n8877), .CK(clk), .Q(reg_mem[940]) );
  DFF_X1 reg_mem_reg_138__3_ ( .D(n8876), .CK(clk), .Q(reg_mem[939]) );
  DFF_X1 reg_mem_reg_138__2_ ( .D(n8875), .CK(clk), .Q(reg_mem[938]) );
  DFF_X1 reg_mem_reg_138__1_ ( .D(n8874), .CK(clk), .Q(reg_mem[937]) );
  DFF_X1 reg_mem_reg_138__0_ ( .D(n8873), .CK(clk), .Q(reg_mem[936]) );
  DFF_X1 reg_mem_reg_139__7_ ( .D(n7151), .CK(clk), .Q(reg_mem[935]) );
  DFF_X1 reg_mem_reg_139__6_ ( .D(n7150), .CK(clk), .Q(reg_mem[934]) );
  DFF_X1 reg_mem_reg_139__5_ ( .D(n7149), .CK(clk), .Q(reg_mem[933]) );
  DFF_X1 reg_mem_reg_139__4_ ( .D(n7148), .CK(clk), .Q(reg_mem[932]) );
  DFF_X1 reg_mem_reg_139__3_ ( .D(n7147), .CK(clk), .Q(reg_mem[931]) );
  DFF_X1 reg_mem_reg_139__2_ ( .D(n7146), .CK(clk), .Q(reg_mem[930]) );
  DFF_X1 reg_mem_reg_139__1_ ( .D(n7145), .CK(clk), .Q(reg_mem[929]) );
  DFF_X1 reg_mem_reg_139__0_ ( .D(n7144), .CK(clk), .Q(reg_mem[928]) );
  DFF_X1 reg_mem_reg_140__7_ ( .D(n8448), .CK(clk), .Q(reg_mem[927]) );
  DFF_X1 reg_mem_reg_140__6_ ( .D(n8447), .CK(clk), .Q(reg_mem[926]) );
  DFF_X1 reg_mem_reg_140__5_ ( .D(n8446), .CK(clk), .Q(reg_mem[925]) );
  DFF_X1 reg_mem_reg_140__4_ ( .D(n8445), .CK(clk), .Q(reg_mem[924]) );
  DFF_X1 reg_mem_reg_140__3_ ( .D(n8444), .CK(clk), .Q(reg_mem[923]) );
  DFF_X1 reg_mem_reg_140__2_ ( .D(n8443), .CK(clk), .Q(reg_mem[922]) );
  DFF_X1 reg_mem_reg_140__1_ ( .D(n8442), .CK(clk), .Q(reg_mem[921]) );
  DFF_X1 reg_mem_reg_140__0_ ( .D(n8441), .CK(clk), .Q(reg_mem[920]) );
  DFF_X1 reg_mem_reg_141__7_ ( .D(n7871), .CK(clk), .Q(reg_mem[919]) );
  DFF_X1 reg_mem_reg_141__6_ ( .D(n7870), .CK(clk), .Q(reg_mem[918]) );
  DFF_X1 reg_mem_reg_141__5_ ( .D(n7869), .CK(clk), .Q(reg_mem[917]) );
  DFF_X1 reg_mem_reg_141__4_ ( .D(n7868), .CK(clk), .Q(reg_mem[916]) );
  DFF_X1 reg_mem_reg_141__3_ ( .D(n7867), .CK(clk), .Q(reg_mem[915]) );
  DFF_X1 reg_mem_reg_141__2_ ( .D(n7866), .CK(clk), .Q(reg_mem[914]) );
  DFF_X1 reg_mem_reg_141__1_ ( .D(n7865), .CK(clk), .Q(reg_mem[913]) );
  DFF_X1 reg_mem_reg_141__0_ ( .D(n7864), .CK(clk), .Q(reg_mem[912]) );
  DFF_X1 reg_mem_reg_142__7_ ( .D(n9024), .CK(clk), .Q(reg_mem[911]) );
  DFF_X1 reg_mem_reg_142__6_ ( .D(n9023), .CK(clk), .Q(reg_mem[910]) );
  DFF_X1 reg_mem_reg_142__5_ ( .D(n9022), .CK(clk), .Q(reg_mem[909]) );
  DFF_X1 reg_mem_reg_142__4_ ( .D(n9021), .CK(clk), .Q(reg_mem[908]) );
  DFF_X1 reg_mem_reg_142__3_ ( .D(n9020), .CK(clk), .Q(reg_mem[907]) );
  DFF_X1 reg_mem_reg_142__2_ ( .D(n9019), .CK(clk), .Q(reg_mem[906]) );
  DFF_X1 reg_mem_reg_142__1_ ( .D(n9018), .CK(clk), .Q(reg_mem[905]) );
  DFF_X1 reg_mem_reg_142__0_ ( .D(n9017), .CK(clk), .Q(reg_mem[904]) );
  DFF_X1 reg_mem_reg_143__7_ ( .D(n7295), .CK(clk), .Q(reg_mem[903]) );
  DFF_X1 reg_mem_reg_143__6_ ( .D(n7294), .CK(clk), .Q(reg_mem[902]) );
  DFF_X1 reg_mem_reg_143__5_ ( .D(n7293), .CK(clk), .Q(reg_mem[901]) );
  DFF_X1 reg_mem_reg_143__4_ ( .D(n7292), .CK(clk), .Q(reg_mem[900]) );
  DFF_X1 reg_mem_reg_143__3_ ( .D(n7291), .CK(clk), .Q(reg_mem[899]) );
  DFF_X1 reg_mem_reg_143__2_ ( .D(n7290), .CK(clk), .Q(reg_mem[898]) );
  DFF_X1 reg_mem_reg_143__1_ ( .D(n7289), .CK(clk), .Q(reg_mem[897]) );
  DFF_X1 reg_mem_reg_143__0_ ( .D(n7288), .CK(clk), .Q(reg_mem[896]) );
  DFF_X1 reg_mem_reg_144__7_ ( .D(n8025), .CK(clk), .Q(reg_mem[895]) );
  DFF_X1 reg_mem_reg_144__6_ ( .D(n8024), .CK(clk), .Q(reg_mem[894]) );
  DFF_X1 reg_mem_reg_144__5_ ( .D(n8023), .CK(clk), .Q(reg_mem[893]) );
  DFF_X1 reg_mem_reg_144__4_ ( .D(n8022), .CK(clk), .Q(reg_mem[892]) );
  DFF_X1 reg_mem_reg_144__3_ ( .D(n8021), .CK(clk), .Q(reg_mem[891]) );
  DFF_X1 reg_mem_reg_144__2_ ( .D(n8020), .CK(clk), .Q(reg_mem[890]) );
  DFF_X1 reg_mem_reg_144__1_ ( .D(n8019), .CK(clk), .Q(reg_mem[889]) );
  DFF_X1 reg_mem_reg_144__0_ ( .D(n8018), .CK(clk), .Q(reg_mem[888]) );
  DFF_X1 reg_mem_reg_145__7_ ( .D(n7448), .CK(clk), .Q(reg_mem[887]) );
  DFF_X1 reg_mem_reg_145__6_ ( .D(n7447), .CK(clk), .Q(reg_mem[886]) );
  DFF_X1 reg_mem_reg_145__5_ ( .D(n7446), .CK(clk), .Q(reg_mem[885]) );
  DFF_X1 reg_mem_reg_145__4_ ( .D(n7445), .CK(clk), .Q(reg_mem[884]) );
  DFF_X1 reg_mem_reg_145__3_ ( .D(n7444), .CK(clk), .Q(reg_mem[883]) );
  DFF_X1 reg_mem_reg_145__2_ ( .D(n7443), .CK(clk), .Q(reg_mem[882]) );
  DFF_X1 reg_mem_reg_145__1_ ( .D(n7442), .CK(clk), .Q(reg_mem[881]) );
  DFF_X1 reg_mem_reg_145__0_ ( .D(n7441), .CK(clk), .Q(reg_mem[880]) );
  DFF_X1 reg_mem_reg_146__7_ ( .D(n8601), .CK(clk), .Q(reg_mem[879]) );
  DFF_X1 reg_mem_reg_146__6_ ( .D(n8600), .CK(clk), .Q(reg_mem[878]) );
  DFF_X1 reg_mem_reg_146__5_ ( .D(n8599), .CK(clk), .Q(reg_mem[877]) );
  DFF_X1 reg_mem_reg_146__4_ ( .D(n8598), .CK(clk), .Q(reg_mem[876]) );
  DFF_X1 reg_mem_reg_146__3_ ( .D(n8597), .CK(clk), .Q(reg_mem[875]) );
  DFF_X1 reg_mem_reg_146__2_ ( .D(n8596), .CK(clk), .Q(reg_mem[874]) );
  DFF_X1 reg_mem_reg_146__1_ ( .D(n8595), .CK(clk), .Q(reg_mem[873]) );
  DFF_X1 reg_mem_reg_146__0_ ( .D(n8594), .CK(clk), .Q(reg_mem[872]) );
  DFF_X1 reg_mem_reg_147__7_ ( .D(n6872), .CK(clk), .Q(reg_mem[871]) );
  DFF_X1 reg_mem_reg_147__6_ ( .D(n6871), .CK(clk), .Q(reg_mem[870]) );
  DFF_X1 reg_mem_reg_147__5_ ( .D(n6870), .CK(clk), .Q(reg_mem[869]) );
  DFF_X1 reg_mem_reg_147__4_ ( .D(n6869), .CK(clk), .Q(reg_mem[868]) );
  DFF_X1 reg_mem_reg_147__3_ ( .D(n6868), .CK(clk), .Q(reg_mem[867]) );
  DFF_X1 reg_mem_reg_147__2_ ( .D(n6867), .CK(clk), .Q(reg_mem[866]) );
  DFF_X1 reg_mem_reg_147__1_ ( .D(n6866), .CK(clk), .Q(reg_mem[865]) );
  DFF_X1 reg_mem_reg_147__0_ ( .D(n6865), .CK(clk), .Q(reg_mem[864]) );
  DFF_X1 reg_mem_reg_148__7_ ( .D(n8169), .CK(clk), .Q(reg_mem[863]) );
  DFF_X1 reg_mem_reg_148__6_ ( .D(n8168), .CK(clk), .Q(reg_mem[862]) );
  DFF_X1 reg_mem_reg_148__5_ ( .D(n8167), .CK(clk), .Q(reg_mem[861]) );
  DFF_X1 reg_mem_reg_148__4_ ( .D(n8166), .CK(clk), .Q(reg_mem[860]) );
  DFF_X1 reg_mem_reg_148__3_ ( .D(n8165), .CK(clk), .Q(reg_mem[859]) );
  DFF_X1 reg_mem_reg_148__2_ ( .D(n8164), .CK(clk), .Q(reg_mem[858]) );
  DFF_X1 reg_mem_reg_148__1_ ( .D(n8163), .CK(clk), .Q(reg_mem[857]) );
  DFF_X1 reg_mem_reg_148__0_ ( .D(n8162), .CK(clk), .Q(reg_mem[856]) );
  DFF_X1 reg_mem_reg_149__7_ ( .D(n7592), .CK(clk), .Q(reg_mem[855]) );
  DFF_X1 reg_mem_reg_149__6_ ( .D(n7591), .CK(clk), .Q(reg_mem[854]) );
  DFF_X1 reg_mem_reg_149__5_ ( .D(n7590), .CK(clk), .Q(reg_mem[853]) );
  DFF_X1 reg_mem_reg_149__4_ ( .D(n7589), .CK(clk), .Q(reg_mem[852]) );
  DFF_X1 reg_mem_reg_149__3_ ( .D(n7588), .CK(clk), .Q(reg_mem[851]) );
  DFF_X1 reg_mem_reg_149__2_ ( .D(n7587), .CK(clk), .Q(reg_mem[850]) );
  DFF_X1 reg_mem_reg_149__1_ ( .D(n7586), .CK(clk), .Q(reg_mem[849]) );
  DFF_X1 reg_mem_reg_149__0_ ( .D(n7585), .CK(clk), .Q(reg_mem[848]) );
  DFF_X1 reg_mem_reg_150__7_ ( .D(n8745), .CK(clk), .Q(reg_mem[847]) );
  DFF_X1 reg_mem_reg_150__6_ ( .D(n8744), .CK(clk), .Q(reg_mem[846]) );
  DFF_X1 reg_mem_reg_150__5_ ( .D(n8743), .CK(clk), .Q(reg_mem[845]) );
  DFF_X1 reg_mem_reg_150__4_ ( .D(n8742), .CK(clk), .Q(reg_mem[844]) );
  DFF_X1 reg_mem_reg_150__3_ ( .D(n8741), .CK(clk), .Q(reg_mem[843]) );
  DFF_X1 reg_mem_reg_150__2_ ( .D(n8740), .CK(clk), .Q(reg_mem[842]) );
  DFF_X1 reg_mem_reg_150__1_ ( .D(n8739), .CK(clk), .Q(reg_mem[841]) );
  DFF_X1 reg_mem_reg_150__0_ ( .D(n8738), .CK(clk), .Q(reg_mem[840]) );
  DFF_X1 reg_mem_reg_151__7_ ( .D(n7016), .CK(clk), .Q(reg_mem[839]) );
  DFF_X1 reg_mem_reg_151__6_ ( .D(n7015), .CK(clk), .Q(reg_mem[838]) );
  DFF_X1 reg_mem_reg_151__5_ ( .D(n7014), .CK(clk), .Q(reg_mem[837]) );
  DFF_X1 reg_mem_reg_151__4_ ( .D(n7013), .CK(clk), .Q(reg_mem[836]) );
  DFF_X1 reg_mem_reg_151__3_ ( .D(n7012), .CK(clk), .Q(reg_mem[835]) );
  DFF_X1 reg_mem_reg_151__2_ ( .D(n7011), .CK(clk), .Q(reg_mem[834]) );
  DFF_X1 reg_mem_reg_151__1_ ( .D(n7010), .CK(clk), .Q(reg_mem[833]) );
  DFF_X1 reg_mem_reg_151__0_ ( .D(n7009), .CK(clk), .Q(reg_mem[832]) );
  DFF_X1 reg_mem_reg_152__7_ ( .D(n8313), .CK(clk), .Q(reg_mem[831]) );
  DFF_X1 reg_mem_reg_152__6_ ( .D(n8312), .CK(clk), .Q(reg_mem[830]) );
  DFF_X1 reg_mem_reg_152__5_ ( .D(n8311), .CK(clk), .Q(reg_mem[829]) );
  DFF_X1 reg_mem_reg_152__4_ ( .D(n8310), .CK(clk), .Q(reg_mem[828]) );
  DFF_X1 reg_mem_reg_152__3_ ( .D(n8309), .CK(clk), .Q(reg_mem[827]) );
  DFF_X1 reg_mem_reg_152__2_ ( .D(n8308), .CK(clk), .Q(reg_mem[826]) );
  DFF_X1 reg_mem_reg_152__1_ ( .D(n8307), .CK(clk), .Q(reg_mem[825]) );
  DFF_X1 reg_mem_reg_152__0_ ( .D(n8306), .CK(clk), .Q(reg_mem[824]) );
  DFF_X1 reg_mem_reg_153__7_ ( .D(n7736), .CK(clk), .Q(reg_mem[823]) );
  DFF_X1 reg_mem_reg_153__6_ ( .D(n7735), .CK(clk), .Q(reg_mem[822]) );
  DFF_X1 reg_mem_reg_153__5_ ( .D(n7734), .CK(clk), .Q(reg_mem[821]) );
  DFF_X1 reg_mem_reg_153__4_ ( .D(n7733), .CK(clk), .Q(reg_mem[820]) );
  DFF_X1 reg_mem_reg_153__3_ ( .D(n7732), .CK(clk), .Q(reg_mem[819]) );
  DFF_X1 reg_mem_reg_153__2_ ( .D(n7731), .CK(clk), .Q(reg_mem[818]) );
  DFF_X1 reg_mem_reg_153__1_ ( .D(n7730), .CK(clk), .Q(reg_mem[817]) );
  DFF_X1 reg_mem_reg_153__0_ ( .D(n7729), .CK(clk), .Q(reg_mem[816]) );
  DFF_X1 reg_mem_reg_154__7_ ( .D(n8889), .CK(clk), .Q(reg_mem[815]) );
  DFF_X1 reg_mem_reg_154__6_ ( .D(n8888), .CK(clk), .Q(reg_mem[814]) );
  DFF_X1 reg_mem_reg_154__5_ ( .D(n8887), .CK(clk), .Q(reg_mem[813]) );
  DFF_X1 reg_mem_reg_154__4_ ( .D(n8886), .CK(clk), .Q(reg_mem[812]) );
  DFF_X1 reg_mem_reg_154__3_ ( .D(n8885), .CK(clk), .Q(reg_mem[811]) );
  DFF_X1 reg_mem_reg_154__2_ ( .D(n8884), .CK(clk), .Q(reg_mem[810]) );
  DFF_X1 reg_mem_reg_154__1_ ( .D(n8883), .CK(clk), .Q(reg_mem[809]) );
  DFF_X1 reg_mem_reg_154__0_ ( .D(n8882), .CK(clk), .Q(reg_mem[808]) );
  DFF_X1 reg_mem_reg_155__7_ ( .D(n7160), .CK(clk), .Q(reg_mem[807]) );
  DFF_X1 reg_mem_reg_155__6_ ( .D(n7159), .CK(clk), .Q(reg_mem[806]) );
  DFF_X1 reg_mem_reg_155__5_ ( .D(n7158), .CK(clk), .Q(reg_mem[805]) );
  DFF_X1 reg_mem_reg_155__4_ ( .D(n7157), .CK(clk), .Q(reg_mem[804]) );
  DFF_X1 reg_mem_reg_155__3_ ( .D(n7156), .CK(clk), .Q(reg_mem[803]) );
  DFF_X1 reg_mem_reg_155__2_ ( .D(n7155), .CK(clk), .Q(reg_mem[802]) );
  DFF_X1 reg_mem_reg_155__1_ ( .D(n7154), .CK(clk), .Q(reg_mem[801]) );
  DFF_X1 reg_mem_reg_155__0_ ( .D(n7153), .CK(clk), .Q(reg_mem[800]) );
  DFF_X1 reg_mem_reg_156__7_ ( .D(n8457), .CK(clk), .Q(reg_mem[799]) );
  DFF_X1 reg_mem_reg_156__6_ ( .D(n8456), .CK(clk), .Q(reg_mem[798]) );
  DFF_X1 reg_mem_reg_156__5_ ( .D(n8455), .CK(clk), .Q(reg_mem[797]) );
  DFF_X1 reg_mem_reg_156__4_ ( .D(n8454), .CK(clk), .Q(reg_mem[796]) );
  DFF_X1 reg_mem_reg_156__3_ ( .D(n8453), .CK(clk), .Q(reg_mem[795]) );
  DFF_X1 reg_mem_reg_156__2_ ( .D(n8452), .CK(clk), .Q(reg_mem[794]) );
  DFF_X1 reg_mem_reg_156__1_ ( .D(n8451), .CK(clk), .Q(reg_mem[793]) );
  DFF_X1 reg_mem_reg_156__0_ ( .D(n8450), .CK(clk), .Q(reg_mem[792]) );
  DFF_X1 reg_mem_reg_157__7_ ( .D(n7880), .CK(clk), .Q(reg_mem[791]) );
  DFF_X1 reg_mem_reg_157__6_ ( .D(n7879), .CK(clk), .Q(reg_mem[790]) );
  DFF_X1 reg_mem_reg_157__5_ ( .D(n7878), .CK(clk), .Q(reg_mem[789]) );
  DFF_X1 reg_mem_reg_157__4_ ( .D(n7877), .CK(clk), .Q(reg_mem[788]) );
  DFF_X1 reg_mem_reg_157__3_ ( .D(n7876), .CK(clk), .Q(reg_mem[787]) );
  DFF_X1 reg_mem_reg_157__2_ ( .D(n7875), .CK(clk), .Q(reg_mem[786]) );
  DFF_X1 reg_mem_reg_157__1_ ( .D(n7874), .CK(clk), .Q(reg_mem[785]) );
  DFF_X1 reg_mem_reg_157__0_ ( .D(n7873), .CK(clk), .Q(reg_mem[784]) );
  DFF_X1 reg_mem_reg_158__7_ ( .D(n9033), .CK(clk), .Q(reg_mem[783]) );
  DFF_X1 reg_mem_reg_158__6_ ( .D(n9032), .CK(clk), .Q(reg_mem[782]) );
  DFF_X1 reg_mem_reg_158__5_ ( .D(n9031), .CK(clk), .Q(reg_mem[781]) );
  DFF_X1 reg_mem_reg_158__4_ ( .D(n9030), .CK(clk), .Q(reg_mem[780]) );
  DFF_X1 reg_mem_reg_158__3_ ( .D(n9029), .CK(clk), .Q(reg_mem[779]) );
  DFF_X1 reg_mem_reg_158__2_ ( .D(n9028), .CK(clk), .Q(reg_mem[778]) );
  DFF_X1 reg_mem_reg_158__1_ ( .D(n9027), .CK(clk), .Q(reg_mem[777]) );
  DFF_X1 reg_mem_reg_158__0_ ( .D(n9026), .CK(clk), .Q(reg_mem[776]) );
  DFF_X1 reg_mem_reg_159__7_ ( .D(n7304), .CK(clk), .Q(reg_mem[775]) );
  DFF_X1 reg_mem_reg_159__6_ ( .D(n7303), .CK(clk), .Q(reg_mem[774]) );
  DFF_X1 reg_mem_reg_159__5_ ( .D(n7302), .CK(clk), .Q(reg_mem[773]) );
  DFF_X1 reg_mem_reg_159__4_ ( .D(n7301), .CK(clk), .Q(reg_mem[772]) );
  DFF_X1 reg_mem_reg_159__3_ ( .D(n7300), .CK(clk), .Q(reg_mem[771]) );
  DFF_X1 reg_mem_reg_159__2_ ( .D(n7299), .CK(clk), .Q(reg_mem[770]) );
  DFF_X1 reg_mem_reg_159__1_ ( .D(n7298), .CK(clk), .Q(reg_mem[769]) );
  DFF_X1 reg_mem_reg_159__0_ ( .D(n7297), .CK(clk), .Q(reg_mem[768]) );
  DFF_X1 reg_mem_reg_160__7_ ( .D(n8034), .CK(clk), .Q(reg_mem[767]) );
  DFF_X1 reg_mem_reg_160__6_ ( .D(n8033), .CK(clk), .Q(reg_mem[766]) );
  DFF_X1 reg_mem_reg_160__5_ ( .D(n8032), .CK(clk), .Q(reg_mem[765]) );
  DFF_X1 reg_mem_reg_160__4_ ( .D(n8031), .CK(clk), .Q(reg_mem[764]) );
  DFF_X1 reg_mem_reg_160__3_ ( .D(n8030), .CK(clk), .Q(reg_mem[763]) );
  DFF_X1 reg_mem_reg_160__2_ ( .D(n8029), .CK(clk), .Q(reg_mem[762]) );
  DFF_X1 reg_mem_reg_160__1_ ( .D(n8028), .CK(clk), .Q(reg_mem[761]) );
  DFF_X1 reg_mem_reg_160__0_ ( .D(n8027), .CK(clk), .Q(reg_mem[760]) );
  DFF_X1 reg_mem_reg_161__7_ ( .D(n7457), .CK(clk), .Q(reg_mem[759]) );
  DFF_X1 reg_mem_reg_161__6_ ( .D(n7456), .CK(clk), .Q(reg_mem[758]) );
  DFF_X1 reg_mem_reg_161__5_ ( .D(n7455), .CK(clk), .Q(reg_mem[757]) );
  DFF_X1 reg_mem_reg_161__4_ ( .D(n7454), .CK(clk), .Q(reg_mem[756]) );
  DFF_X1 reg_mem_reg_161__3_ ( .D(n7453), .CK(clk), .Q(reg_mem[755]) );
  DFF_X1 reg_mem_reg_161__2_ ( .D(n7452), .CK(clk), .Q(reg_mem[754]) );
  DFF_X1 reg_mem_reg_161__1_ ( .D(n7451), .CK(clk), .Q(reg_mem[753]) );
  DFF_X1 reg_mem_reg_161__0_ ( .D(n7450), .CK(clk), .Q(reg_mem[752]) );
  DFF_X1 reg_mem_reg_162__7_ ( .D(n8610), .CK(clk), .Q(reg_mem[751]) );
  DFF_X1 reg_mem_reg_162__6_ ( .D(n8609), .CK(clk), .Q(reg_mem[750]) );
  DFF_X1 reg_mem_reg_162__5_ ( .D(n8608), .CK(clk), .Q(reg_mem[749]) );
  DFF_X1 reg_mem_reg_162__4_ ( .D(n8607), .CK(clk), .Q(reg_mem[748]) );
  DFF_X1 reg_mem_reg_162__3_ ( .D(n8606), .CK(clk), .Q(reg_mem[747]) );
  DFF_X1 reg_mem_reg_162__2_ ( .D(n8605), .CK(clk), .Q(reg_mem[746]) );
  DFF_X1 reg_mem_reg_162__1_ ( .D(n8604), .CK(clk), .Q(reg_mem[745]) );
  DFF_X1 reg_mem_reg_162__0_ ( .D(n8603), .CK(clk), .Q(reg_mem[744]) );
  DFF_X1 reg_mem_reg_163__7_ ( .D(n6881), .CK(clk), .Q(reg_mem[743]) );
  DFF_X1 reg_mem_reg_163__6_ ( .D(n6880), .CK(clk), .Q(reg_mem[742]) );
  DFF_X1 reg_mem_reg_163__5_ ( .D(n6879), .CK(clk), .Q(reg_mem[741]) );
  DFF_X1 reg_mem_reg_163__4_ ( .D(n6878), .CK(clk), .Q(reg_mem[740]) );
  DFF_X1 reg_mem_reg_163__3_ ( .D(n6877), .CK(clk), .Q(reg_mem[739]) );
  DFF_X1 reg_mem_reg_163__2_ ( .D(n6876), .CK(clk), .Q(reg_mem[738]) );
  DFF_X1 reg_mem_reg_163__1_ ( .D(n6875), .CK(clk), .Q(reg_mem[737]) );
  DFF_X1 reg_mem_reg_163__0_ ( .D(n6874), .CK(clk), .Q(reg_mem[736]) );
  DFF_X1 reg_mem_reg_164__7_ ( .D(n8178), .CK(clk), .Q(reg_mem[735]) );
  DFF_X1 reg_mem_reg_164__6_ ( .D(n8177), .CK(clk), .Q(reg_mem[734]) );
  DFF_X1 reg_mem_reg_164__5_ ( .D(n8176), .CK(clk), .Q(reg_mem[733]) );
  DFF_X1 reg_mem_reg_164__4_ ( .D(n8175), .CK(clk), .Q(reg_mem[732]) );
  DFF_X1 reg_mem_reg_164__3_ ( .D(n8174), .CK(clk), .Q(reg_mem[731]) );
  DFF_X1 reg_mem_reg_164__2_ ( .D(n8173), .CK(clk), .Q(reg_mem[730]) );
  DFF_X1 reg_mem_reg_164__1_ ( .D(n8172), .CK(clk), .Q(reg_mem[729]) );
  DFF_X1 reg_mem_reg_164__0_ ( .D(n8171), .CK(clk), .Q(reg_mem[728]) );
  DFF_X1 reg_mem_reg_165__7_ ( .D(n7601), .CK(clk), .Q(reg_mem[727]) );
  DFF_X1 reg_mem_reg_165__6_ ( .D(n7600), .CK(clk), .Q(reg_mem[726]) );
  DFF_X1 reg_mem_reg_165__5_ ( .D(n7599), .CK(clk), .Q(reg_mem[725]) );
  DFF_X1 reg_mem_reg_165__4_ ( .D(n7598), .CK(clk), .Q(reg_mem[724]) );
  DFF_X1 reg_mem_reg_165__3_ ( .D(n7597), .CK(clk), .Q(reg_mem[723]) );
  DFF_X1 reg_mem_reg_165__2_ ( .D(n7596), .CK(clk), .Q(reg_mem[722]) );
  DFF_X1 reg_mem_reg_165__1_ ( .D(n7595), .CK(clk), .Q(reg_mem[721]) );
  DFF_X1 reg_mem_reg_165__0_ ( .D(n7594), .CK(clk), .Q(reg_mem[720]) );
  DFF_X1 reg_mem_reg_166__7_ ( .D(n8754), .CK(clk), .Q(reg_mem[719]) );
  DFF_X1 reg_mem_reg_166__6_ ( .D(n8753), .CK(clk), .Q(reg_mem[718]) );
  DFF_X1 reg_mem_reg_166__5_ ( .D(n8752), .CK(clk), .Q(reg_mem[717]) );
  DFF_X1 reg_mem_reg_166__4_ ( .D(n8751), .CK(clk), .Q(reg_mem[716]) );
  DFF_X1 reg_mem_reg_166__3_ ( .D(n8750), .CK(clk), .Q(reg_mem[715]) );
  DFF_X1 reg_mem_reg_166__2_ ( .D(n8749), .CK(clk), .Q(reg_mem[714]) );
  DFF_X1 reg_mem_reg_166__1_ ( .D(n8748), .CK(clk), .Q(reg_mem[713]) );
  DFF_X1 reg_mem_reg_166__0_ ( .D(n8747), .CK(clk), .Q(reg_mem[712]) );
  DFF_X1 reg_mem_reg_167__7_ ( .D(n7025), .CK(clk), .Q(reg_mem[711]) );
  DFF_X1 reg_mem_reg_167__6_ ( .D(n7024), .CK(clk), .Q(reg_mem[710]) );
  DFF_X1 reg_mem_reg_167__5_ ( .D(n7023), .CK(clk), .Q(reg_mem[709]) );
  DFF_X1 reg_mem_reg_167__4_ ( .D(n7022), .CK(clk), .Q(reg_mem[708]) );
  DFF_X1 reg_mem_reg_167__3_ ( .D(n7021), .CK(clk), .Q(reg_mem[707]) );
  DFF_X1 reg_mem_reg_167__2_ ( .D(n7020), .CK(clk), .Q(reg_mem[706]) );
  DFF_X1 reg_mem_reg_167__1_ ( .D(n7019), .CK(clk), .Q(reg_mem[705]) );
  DFF_X1 reg_mem_reg_167__0_ ( .D(n7018), .CK(clk), .Q(reg_mem[704]) );
  DFF_X1 reg_mem_reg_168__7_ ( .D(n8322), .CK(clk), .Q(reg_mem[703]) );
  DFF_X1 reg_mem_reg_168__6_ ( .D(n8321), .CK(clk), .Q(reg_mem[702]) );
  DFF_X1 reg_mem_reg_168__5_ ( .D(n8320), .CK(clk), .Q(reg_mem[701]) );
  DFF_X1 reg_mem_reg_168__4_ ( .D(n8319), .CK(clk), .Q(reg_mem[700]) );
  DFF_X1 reg_mem_reg_168__3_ ( .D(n8318), .CK(clk), .Q(reg_mem[699]) );
  DFF_X1 reg_mem_reg_168__2_ ( .D(n8317), .CK(clk), .Q(reg_mem[698]) );
  DFF_X1 reg_mem_reg_168__1_ ( .D(n8316), .CK(clk), .Q(reg_mem[697]) );
  DFF_X1 reg_mem_reg_168__0_ ( .D(n8315), .CK(clk), .Q(reg_mem[696]) );
  DFF_X1 reg_mem_reg_169__7_ ( .D(n7745), .CK(clk), .Q(reg_mem[695]) );
  DFF_X1 reg_mem_reg_169__6_ ( .D(n7744), .CK(clk), .Q(reg_mem[694]) );
  DFF_X1 reg_mem_reg_169__5_ ( .D(n7743), .CK(clk), .Q(reg_mem[693]) );
  DFF_X1 reg_mem_reg_169__4_ ( .D(n7742), .CK(clk), .Q(reg_mem[692]) );
  DFF_X1 reg_mem_reg_169__3_ ( .D(n7741), .CK(clk), .Q(reg_mem[691]) );
  DFF_X1 reg_mem_reg_169__2_ ( .D(n7740), .CK(clk), .Q(reg_mem[690]) );
  DFF_X1 reg_mem_reg_169__1_ ( .D(n7739), .CK(clk), .Q(reg_mem[689]) );
  DFF_X1 reg_mem_reg_169__0_ ( .D(n7738), .CK(clk), .Q(reg_mem[688]) );
  DFF_X1 reg_mem_reg_170__7_ ( .D(n8898), .CK(clk), .Q(reg_mem[687]) );
  DFF_X1 reg_mem_reg_170__6_ ( .D(n8897), .CK(clk), .Q(reg_mem[686]) );
  DFF_X1 reg_mem_reg_170__5_ ( .D(n8896), .CK(clk), .Q(reg_mem[685]) );
  DFF_X1 reg_mem_reg_170__4_ ( .D(n8895), .CK(clk), .Q(reg_mem[684]) );
  DFF_X1 reg_mem_reg_170__3_ ( .D(n8894), .CK(clk), .Q(reg_mem[683]) );
  DFF_X1 reg_mem_reg_170__2_ ( .D(n8893), .CK(clk), .Q(reg_mem[682]) );
  DFF_X1 reg_mem_reg_170__1_ ( .D(n8892), .CK(clk), .Q(reg_mem[681]) );
  DFF_X1 reg_mem_reg_170__0_ ( .D(n8891), .CK(clk), .Q(reg_mem[680]) );
  DFF_X1 reg_mem_reg_171__7_ ( .D(n7169), .CK(clk), .Q(reg_mem[679]) );
  DFF_X1 reg_mem_reg_171__6_ ( .D(n7168), .CK(clk), .Q(reg_mem[678]) );
  DFF_X1 reg_mem_reg_171__5_ ( .D(n7167), .CK(clk), .Q(reg_mem[677]) );
  DFF_X1 reg_mem_reg_171__4_ ( .D(n7166), .CK(clk), .Q(reg_mem[676]) );
  DFF_X1 reg_mem_reg_171__3_ ( .D(n7165), .CK(clk), .Q(reg_mem[675]) );
  DFF_X1 reg_mem_reg_171__2_ ( .D(n7164), .CK(clk), .Q(reg_mem[674]) );
  DFF_X1 reg_mem_reg_171__1_ ( .D(n7163), .CK(clk), .Q(reg_mem[673]) );
  DFF_X1 reg_mem_reg_171__0_ ( .D(n7162), .CK(clk), .Q(reg_mem[672]) );
  DFF_X1 reg_mem_reg_172__7_ ( .D(n8466), .CK(clk), .Q(reg_mem[671]) );
  DFF_X1 reg_mem_reg_172__6_ ( .D(n8465), .CK(clk), .Q(reg_mem[670]) );
  DFF_X1 reg_mem_reg_172__5_ ( .D(n8464), .CK(clk), .Q(reg_mem[669]) );
  DFF_X1 reg_mem_reg_172__4_ ( .D(n8463), .CK(clk), .Q(reg_mem[668]) );
  DFF_X1 reg_mem_reg_172__3_ ( .D(n8462), .CK(clk), .Q(reg_mem[667]) );
  DFF_X1 reg_mem_reg_172__2_ ( .D(n8461), .CK(clk), .Q(reg_mem[666]) );
  DFF_X1 reg_mem_reg_172__1_ ( .D(n8460), .CK(clk), .Q(reg_mem[665]) );
  DFF_X1 reg_mem_reg_172__0_ ( .D(n8459), .CK(clk), .Q(reg_mem[664]) );
  DFF_X1 reg_mem_reg_173__7_ ( .D(n7889), .CK(clk), .Q(reg_mem[663]) );
  DFF_X1 reg_mem_reg_173__6_ ( .D(n7888), .CK(clk), .Q(reg_mem[662]) );
  DFF_X1 reg_mem_reg_173__5_ ( .D(n7887), .CK(clk), .Q(reg_mem[661]) );
  DFF_X1 reg_mem_reg_173__4_ ( .D(n7886), .CK(clk), .Q(reg_mem[660]) );
  DFF_X1 reg_mem_reg_173__3_ ( .D(n7885), .CK(clk), .Q(reg_mem[659]) );
  DFF_X1 reg_mem_reg_173__2_ ( .D(n7884), .CK(clk), .Q(reg_mem[658]) );
  DFF_X1 reg_mem_reg_173__1_ ( .D(n7883), .CK(clk), .Q(reg_mem[657]) );
  DFF_X1 reg_mem_reg_173__0_ ( .D(n7882), .CK(clk), .Q(reg_mem[656]) );
  DFF_X1 reg_mem_reg_174__7_ ( .D(n9042), .CK(clk), .Q(reg_mem[655]) );
  DFF_X1 reg_mem_reg_174__6_ ( .D(n9041), .CK(clk), .Q(reg_mem[654]) );
  DFF_X1 reg_mem_reg_174__5_ ( .D(n9040), .CK(clk), .Q(reg_mem[653]) );
  DFF_X1 reg_mem_reg_174__4_ ( .D(n9039), .CK(clk), .Q(reg_mem[652]) );
  DFF_X1 reg_mem_reg_174__3_ ( .D(n9038), .CK(clk), .Q(reg_mem[651]) );
  DFF_X1 reg_mem_reg_174__2_ ( .D(n9037), .CK(clk), .Q(reg_mem[650]) );
  DFF_X1 reg_mem_reg_174__1_ ( .D(n9036), .CK(clk), .Q(reg_mem[649]) );
  DFF_X1 reg_mem_reg_174__0_ ( .D(n9035), .CK(clk), .Q(reg_mem[648]) );
  DFF_X1 reg_mem_reg_175__7_ ( .D(n7313), .CK(clk), .Q(reg_mem[647]) );
  DFF_X1 reg_mem_reg_175__6_ ( .D(n7312), .CK(clk), .Q(reg_mem[646]) );
  DFF_X1 reg_mem_reg_175__5_ ( .D(n7311), .CK(clk), .Q(reg_mem[645]) );
  DFF_X1 reg_mem_reg_175__4_ ( .D(n7310), .CK(clk), .Q(reg_mem[644]) );
  DFF_X1 reg_mem_reg_175__3_ ( .D(n7309), .CK(clk), .Q(reg_mem[643]) );
  DFF_X1 reg_mem_reg_175__2_ ( .D(n7308), .CK(clk), .Q(reg_mem[642]) );
  DFF_X1 reg_mem_reg_175__1_ ( .D(n7307), .CK(clk), .Q(reg_mem[641]) );
  DFF_X1 reg_mem_reg_175__0_ ( .D(n7306), .CK(clk), .Q(reg_mem[640]) );
  DFF_X1 reg_mem_reg_176__7_ ( .D(n8043), .CK(clk), .Q(reg_mem[639]) );
  DFF_X1 reg_mem_reg_176__6_ ( .D(n8042), .CK(clk), .Q(reg_mem[638]) );
  DFF_X1 reg_mem_reg_176__5_ ( .D(n8041), .CK(clk), .Q(reg_mem[637]) );
  DFF_X1 reg_mem_reg_176__4_ ( .D(n8040), .CK(clk), .Q(reg_mem[636]) );
  DFF_X1 reg_mem_reg_176__3_ ( .D(n8039), .CK(clk), .Q(reg_mem[635]) );
  DFF_X1 reg_mem_reg_176__2_ ( .D(n8038), .CK(clk), .Q(reg_mem[634]) );
  DFF_X1 reg_mem_reg_176__1_ ( .D(n8037), .CK(clk), .Q(reg_mem[633]) );
  DFF_X1 reg_mem_reg_176__0_ ( .D(n8036), .CK(clk), .Q(reg_mem[632]) );
  DFF_X1 reg_mem_reg_177__7_ ( .D(n7466), .CK(clk), .Q(reg_mem[631]) );
  DFF_X1 reg_mem_reg_177__6_ ( .D(n7465), .CK(clk), .Q(reg_mem[630]) );
  DFF_X1 reg_mem_reg_177__5_ ( .D(n7464), .CK(clk), .Q(reg_mem[629]) );
  DFF_X1 reg_mem_reg_177__4_ ( .D(n7463), .CK(clk), .Q(reg_mem[628]) );
  DFF_X1 reg_mem_reg_177__3_ ( .D(n7462), .CK(clk), .Q(reg_mem[627]) );
  DFF_X1 reg_mem_reg_177__2_ ( .D(n7461), .CK(clk), .Q(reg_mem[626]) );
  DFF_X1 reg_mem_reg_177__1_ ( .D(n7460), .CK(clk), .Q(reg_mem[625]) );
  DFF_X1 reg_mem_reg_177__0_ ( .D(n7459), .CK(clk), .Q(reg_mem[624]) );
  DFF_X1 reg_mem_reg_178__7_ ( .D(n8619), .CK(clk), .Q(reg_mem[623]) );
  DFF_X1 reg_mem_reg_178__6_ ( .D(n8618), .CK(clk), .Q(reg_mem[622]) );
  DFF_X1 reg_mem_reg_178__5_ ( .D(n8617), .CK(clk), .Q(reg_mem[621]) );
  DFF_X1 reg_mem_reg_178__4_ ( .D(n8616), .CK(clk), .Q(reg_mem[620]) );
  DFF_X1 reg_mem_reg_178__3_ ( .D(n8615), .CK(clk), .Q(reg_mem[619]) );
  DFF_X1 reg_mem_reg_178__2_ ( .D(n8614), .CK(clk), .Q(reg_mem[618]) );
  DFF_X1 reg_mem_reg_178__1_ ( .D(n8613), .CK(clk), .Q(reg_mem[617]) );
  DFF_X1 reg_mem_reg_178__0_ ( .D(n8612), .CK(clk), .Q(reg_mem[616]) );
  DFF_X1 reg_mem_reg_179__7_ ( .D(n6890), .CK(clk), .Q(reg_mem[615]) );
  DFF_X1 reg_mem_reg_179__6_ ( .D(n6889), .CK(clk), .Q(reg_mem[614]) );
  DFF_X1 reg_mem_reg_179__5_ ( .D(n6888), .CK(clk), .Q(reg_mem[613]) );
  DFF_X1 reg_mem_reg_179__4_ ( .D(n6887), .CK(clk), .Q(reg_mem[612]) );
  DFF_X1 reg_mem_reg_179__3_ ( .D(n6886), .CK(clk), .Q(reg_mem[611]) );
  DFF_X1 reg_mem_reg_179__2_ ( .D(n6885), .CK(clk), .Q(reg_mem[610]) );
  DFF_X1 reg_mem_reg_179__1_ ( .D(n6884), .CK(clk), .Q(reg_mem[609]) );
  DFF_X1 reg_mem_reg_179__0_ ( .D(n6883), .CK(clk), .Q(reg_mem[608]) );
  DFF_X1 reg_mem_reg_180__7_ ( .D(n8187), .CK(clk), .Q(reg_mem[607]) );
  DFF_X1 reg_mem_reg_180__6_ ( .D(n8186), .CK(clk), .Q(reg_mem[606]) );
  DFF_X1 reg_mem_reg_180__5_ ( .D(n8185), .CK(clk), .Q(reg_mem[605]) );
  DFF_X1 reg_mem_reg_180__4_ ( .D(n8184), .CK(clk), .Q(reg_mem[604]) );
  DFF_X1 reg_mem_reg_180__3_ ( .D(n8183), .CK(clk), .Q(reg_mem[603]) );
  DFF_X1 reg_mem_reg_180__2_ ( .D(n8182), .CK(clk), .Q(reg_mem[602]) );
  DFF_X1 reg_mem_reg_180__1_ ( .D(n8181), .CK(clk), .Q(reg_mem[601]) );
  DFF_X1 reg_mem_reg_180__0_ ( .D(n8180), .CK(clk), .Q(reg_mem[600]) );
  DFF_X1 reg_mem_reg_181__7_ ( .D(n7610), .CK(clk), .Q(reg_mem[599]) );
  DFF_X1 reg_mem_reg_181__6_ ( .D(n7609), .CK(clk), .Q(reg_mem[598]) );
  DFF_X1 reg_mem_reg_181__5_ ( .D(n7608), .CK(clk), .Q(reg_mem[597]) );
  DFF_X1 reg_mem_reg_181__4_ ( .D(n7607), .CK(clk), .Q(reg_mem[596]) );
  DFF_X1 reg_mem_reg_181__3_ ( .D(n7606), .CK(clk), .Q(reg_mem[595]) );
  DFF_X1 reg_mem_reg_181__2_ ( .D(n7605), .CK(clk), .Q(reg_mem[594]) );
  DFF_X1 reg_mem_reg_181__1_ ( .D(n7604), .CK(clk), .Q(reg_mem[593]) );
  DFF_X1 reg_mem_reg_181__0_ ( .D(n7603), .CK(clk), .Q(reg_mem[592]) );
  DFF_X1 reg_mem_reg_182__7_ ( .D(n8763), .CK(clk), .Q(reg_mem[591]) );
  DFF_X1 reg_mem_reg_182__6_ ( .D(n8762), .CK(clk), .Q(reg_mem[590]) );
  DFF_X1 reg_mem_reg_182__5_ ( .D(n8761), .CK(clk), .Q(reg_mem[589]) );
  DFF_X1 reg_mem_reg_182__4_ ( .D(n8760), .CK(clk), .Q(reg_mem[588]) );
  DFF_X1 reg_mem_reg_182__3_ ( .D(n8759), .CK(clk), .Q(reg_mem[587]) );
  DFF_X1 reg_mem_reg_182__2_ ( .D(n8758), .CK(clk), .Q(reg_mem[586]) );
  DFF_X1 reg_mem_reg_182__1_ ( .D(n8757), .CK(clk), .Q(reg_mem[585]) );
  DFF_X1 reg_mem_reg_182__0_ ( .D(n8756), .CK(clk), .Q(reg_mem[584]) );
  DFF_X1 reg_mem_reg_183__7_ ( .D(n7034), .CK(clk), .Q(reg_mem[583]) );
  DFF_X1 reg_mem_reg_183__6_ ( .D(n7033), .CK(clk), .Q(reg_mem[582]) );
  DFF_X1 reg_mem_reg_183__5_ ( .D(n7032), .CK(clk), .Q(reg_mem[581]) );
  DFF_X1 reg_mem_reg_183__4_ ( .D(n7031), .CK(clk), .Q(reg_mem[580]) );
  DFF_X1 reg_mem_reg_183__3_ ( .D(n7030), .CK(clk), .Q(reg_mem[579]) );
  DFF_X1 reg_mem_reg_183__2_ ( .D(n7029), .CK(clk), .Q(reg_mem[578]) );
  DFF_X1 reg_mem_reg_183__1_ ( .D(n7028), .CK(clk), .Q(reg_mem[577]) );
  DFF_X1 reg_mem_reg_183__0_ ( .D(n7027), .CK(clk), .Q(reg_mem[576]) );
  DFF_X1 reg_mem_reg_184__7_ ( .D(n8331), .CK(clk), .Q(reg_mem[575]) );
  DFF_X1 reg_mem_reg_184__6_ ( .D(n8330), .CK(clk), .Q(reg_mem[574]) );
  DFF_X1 reg_mem_reg_184__5_ ( .D(n8329), .CK(clk), .Q(reg_mem[573]) );
  DFF_X1 reg_mem_reg_184__4_ ( .D(n8328), .CK(clk), .Q(reg_mem[572]) );
  DFF_X1 reg_mem_reg_184__3_ ( .D(n8327), .CK(clk), .Q(reg_mem[571]) );
  DFF_X1 reg_mem_reg_184__2_ ( .D(n8326), .CK(clk), .Q(reg_mem[570]) );
  DFF_X1 reg_mem_reg_184__1_ ( .D(n8325), .CK(clk), .Q(reg_mem[569]) );
  DFF_X1 reg_mem_reg_184__0_ ( .D(n8324), .CK(clk), .Q(reg_mem[568]) );
  DFF_X1 reg_mem_reg_185__7_ ( .D(n7754), .CK(clk), .Q(reg_mem[567]) );
  DFF_X1 reg_mem_reg_185__6_ ( .D(n7753), .CK(clk), .Q(reg_mem[566]) );
  DFF_X1 reg_mem_reg_185__5_ ( .D(n7752), .CK(clk), .Q(reg_mem[565]) );
  DFF_X1 reg_mem_reg_185__4_ ( .D(n7751), .CK(clk), .Q(reg_mem[564]) );
  DFF_X1 reg_mem_reg_185__3_ ( .D(n7750), .CK(clk), .Q(reg_mem[563]) );
  DFF_X1 reg_mem_reg_185__2_ ( .D(n7749), .CK(clk), .Q(reg_mem[562]) );
  DFF_X1 reg_mem_reg_185__1_ ( .D(n7748), .CK(clk), .Q(reg_mem[561]) );
  DFF_X1 reg_mem_reg_185__0_ ( .D(n7747), .CK(clk), .Q(reg_mem[560]) );
  DFF_X1 reg_mem_reg_186__7_ ( .D(n8907), .CK(clk), .Q(reg_mem[559]) );
  DFF_X1 reg_mem_reg_186__6_ ( .D(n8906), .CK(clk), .Q(reg_mem[558]) );
  DFF_X1 reg_mem_reg_186__5_ ( .D(n8905), .CK(clk), .Q(reg_mem[557]) );
  DFF_X1 reg_mem_reg_186__4_ ( .D(n8904), .CK(clk), .Q(reg_mem[556]) );
  DFF_X1 reg_mem_reg_186__3_ ( .D(n8903), .CK(clk), .Q(reg_mem[555]) );
  DFF_X1 reg_mem_reg_186__2_ ( .D(n8902), .CK(clk), .Q(reg_mem[554]) );
  DFF_X1 reg_mem_reg_186__1_ ( .D(n8901), .CK(clk), .Q(reg_mem[553]) );
  DFF_X1 reg_mem_reg_186__0_ ( .D(n8900), .CK(clk), .Q(reg_mem[552]) );
  DFF_X1 reg_mem_reg_187__7_ ( .D(n7178), .CK(clk), .Q(reg_mem[551]) );
  DFF_X1 reg_mem_reg_187__6_ ( .D(n7177), .CK(clk), .Q(reg_mem[550]) );
  DFF_X1 reg_mem_reg_187__5_ ( .D(n7176), .CK(clk), .Q(reg_mem[549]) );
  DFF_X1 reg_mem_reg_187__4_ ( .D(n7175), .CK(clk), .Q(reg_mem[548]) );
  DFF_X1 reg_mem_reg_187__3_ ( .D(n7174), .CK(clk), .Q(reg_mem[547]) );
  DFF_X1 reg_mem_reg_187__2_ ( .D(n7173), .CK(clk), .Q(reg_mem[546]) );
  DFF_X1 reg_mem_reg_187__1_ ( .D(n7172), .CK(clk), .Q(reg_mem[545]) );
  DFF_X1 reg_mem_reg_187__0_ ( .D(n7171), .CK(clk), .Q(reg_mem[544]) );
  DFF_X1 reg_mem_reg_188__7_ ( .D(n8475), .CK(clk), .Q(reg_mem[543]) );
  DFF_X1 reg_mem_reg_188__6_ ( .D(n8474), .CK(clk), .Q(reg_mem[542]) );
  DFF_X1 reg_mem_reg_188__5_ ( .D(n8473), .CK(clk), .Q(reg_mem[541]) );
  DFF_X1 reg_mem_reg_188__4_ ( .D(n8472), .CK(clk), .Q(reg_mem[540]) );
  DFF_X1 reg_mem_reg_188__3_ ( .D(n8471), .CK(clk), .Q(reg_mem[539]) );
  DFF_X1 reg_mem_reg_188__2_ ( .D(n8470), .CK(clk), .Q(reg_mem[538]) );
  DFF_X1 reg_mem_reg_188__1_ ( .D(n8469), .CK(clk), .Q(reg_mem[537]) );
  DFF_X1 reg_mem_reg_188__0_ ( .D(n8468), .CK(clk), .Q(reg_mem[536]) );
  DFF_X1 reg_mem_reg_189__7_ ( .D(n7898), .CK(clk), .Q(reg_mem[535]) );
  DFF_X1 reg_mem_reg_189__6_ ( .D(n7897), .CK(clk), .Q(reg_mem[534]) );
  DFF_X1 reg_mem_reg_189__5_ ( .D(n7896), .CK(clk), .Q(reg_mem[533]) );
  DFF_X1 reg_mem_reg_189__4_ ( .D(n7895), .CK(clk), .Q(reg_mem[532]) );
  DFF_X1 reg_mem_reg_189__3_ ( .D(n7894), .CK(clk), .Q(reg_mem[531]) );
  DFF_X1 reg_mem_reg_189__2_ ( .D(n7893), .CK(clk), .Q(reg_mem[530]) );
  DFF_X1 reg_mem_reg_189__1_ ( .D(n7892), .CK(clk), .Q(reg_mem[529]) );
  DFF_X1 reg_mem_reg_189__0_ ( .D(n7891), .CK(clk), .Q(reg_mem[528]) );
  DFF_X1 reg_mem_reg_190__7_ ( .D(n9051), .CK(clk), .Q(reg_mem[527]) );
  DFF_X1 reg_mem_reg_190__6_ ( .D(n9050), .CK(clk), .Q(reg_mem[526]) );
  DFF_X1 reg_mem_reg_190__5_ ( .D(n9049), .CK(clk), .Q(reg_mem[525]) );
  DFF_X1 reg_mem_reg_190__4_ ( .D(n9048), .CK(clk), .Q(reg_mem[524]) );
  DFF_X1 reg_mem_reg_190__3_ ( .D(n9047), .CK(clk), .Q(reg_mem[523]) );
  DFF_X1 reg_mem_reg_190__2_ ( .D(n9046), .CK(clk), .Q(reg_mem[522]) );
  DFF_X1 reg_mem_reg_190__1_ ( .D(n9045), .CK(clk), .Q(reg_mem[521]) );
  DFF_X1 reg_mem_reg_190__0_ ( .D(n9044), .CK(clk), .Q(reg_mem[520]) );
  DFF_X1 reg_mem_reg_191__7_ ( .D(n7322), .CK(clk), .Q(reg_mem[519]) );
  DFF_X1 reg_mem_reg_191__6_ ( .D(n7321), .CK(clk), .Q(reg_mem[518]) );
  DFF_X1 reg_mem_reg_191__5_ ( .D(n7320), .CK(clk), .Q(reg_mem[517]) );
  DFF_X1 reg_mem_reg_191__4_ ( .D(n7319), .CK(clk), .Q(reg_mem[516]) );
  DFF_X1 reg_mem_reg_191__3_ ( .D(n7318), .CK(clk), .Q(reg_mem[515]) );
  DFF_X1 reg_mem_reg_191__2_ ( .D(n7317), .CK(clk), .Q(reg_mem[514]) );
  DFF_X1 reg_mem_reg_191__1_ ( .D(n7316), .CK(clk), .Q(reg_mem[513]) );
  DFF_X1 reg_mem_reg_191__0_ ( .D(n7315), .CK(clk), .Q(reg_mem[512]) );
  DFF_X1 reg_mem_reg_192__7_ ( .D(n8052), .CK(clk), .Q(reg_mem[511]) );
  DFF_X1 reg_mem_reg_192__6_ ( .D(n8051), .CK(clk), .Q(reg_mem[510]) );
  DFF_X1 reg_mem_reg_192__5_ ( .D(n8050), .CK(clk), .Q(reg_mem[509]) );
  DFF_X1 reg_mem_reg_192__4_ ( .D(n8049), .CK(clk), .Q(reg_mem[508]) );
  DFF_X1 reg_mem_reg_192__3_ ( .D(n8048), .CK(clk), .Q(reg_mem[507]) );
  DFF_X1 reg_mem_reg_192__2_ ( .D(n8047), .CK(clk), .Q(reg_mem[506]) );
  DFF_X1 reg_mem_reg_192__1_ ( .D(n8046), .CK(clk), .Q(reg_mem[505]) );
  DFF_X1 reg_mem_reg_192__0_ ( .D(n8045), .CK(clk), .Q(reg_mem[504]) );
  DFF_X1 reg_mem_reg_193__7_ ( .D(n7475), .CK(clk), .Q(reg_mem[503]) );
  DFF_X1 reg_mem_reg_193__6_ ( .D(n7474), .CK(clk), .Q(reg_mem[502]) );
  DFF_X1 reg_mem_reg_193__5_ ( .D(n7473), .CK(clk), .Q(reg_mem[501]) );
  DFF_X1 reg_mem_reg_193__4_ ( .D(n7472), .CK(clk), .Q(reg_mem[500]) );
  DFF_X1 reg_mem_reg_193__3_ ( .D(n7471), .CK(clk), .Q(reg_mem[499]) );
  DFF_X1 reg_mem_reg_193__2_ ( .D(n7470), .CK(clk), .Q(reg_mem[498]) );
  DFF_X1 reg_mem_reg_193__1_ ( .D(n7469), .CK(clk), .Q(reg_mem[497]) );
  DFF_X1 reg_mem_reg_193__0_ ( .D(n7468), .CK(clk), .Q(reg_mem[496]) );
  DFF_X1 reg_mem_reg_194__7_ ( .D(n8628), .CK(clk), .Q(reg_mem[495]) );
  DFF_X1 reg_mem_reg_194__6_ ( .D(n8627), .CK(clk), .Q(reg_mem[494]) );
  DFF_X1 reg_mem_reg_194__5_ ( .D(n8626), .CK(clk), .Q(reg_mem[493]) );
  DFF_X1 reg_mem_reg_194__4_ ( .D(n8625), .CK(clk), .Q(reg_mem[492]) );
  DFF_X1 reg_mem_reg_194__3_ ( .D(n8624), .CK(clk), .Q(reg_mem[491]) );
  DFF_X1 reg_mem_reg_194__2_ ( .D(n8623), .CK(clk), .Q(reg_mem[490]) );
  DFF_X1 reg_mem_reg_194__1_ ( .D(n8622), .CK(clk), .Q(reg_mem[489]) );
  DFF_X1 reg_mem_reg_194__0_ ( .D(n8621), .CK(clk), .Q(reg_mem[488]) );
  DFF_X1 reg_mem_reg_195__7_ ( .D(n6899), .CK(clk), .Q(reg_mem[487]) );
  DFF_X1 reg_mem_reg_195__6_ ( .D(n6898), .CK(clk), .Q(reg_mem[486]) );
  DFF_X1 reg_mem_reg_195__5_ ( .D(n6897), .CK(clk), .Q(reg_mem[485]) );
  DFF_X1 reg_mem_reg_195__4_ ( .D(n6896), .CK(clk), .Q(reg_mem[484]) );
  DFF_X1 reg_mem_reg_195__3_ ( .D(n6895), .CK(clk), .Q(reg_mem[483]) );
  DFF_X1 reg_mem_reg_195__2_ ( .D(n6894), .CK(clk), .Q(reg_mem[482]) );
  DFF_X1 reg_mem_reg_195__1_ ( .D(n6893), .CK(clk), .Q(reg_mem[481]) );
  DFF_X1 reg_mem_reg_195__0_ ( .D(n6892), .CK(clk), .Q(reg_mem[480]) );
  DFF_X1 reg_mem_reg_196__7_ ( .D(n8196), .CK(clk), .Q(reg_mem[479]) );
  DFF_X1 reg_mem_reg_196__6_ ( .D(n8195), .CK(clk), .Q(reg_mem[478]) );
  DFF_X1 reg_mem_reg_196__5_ ( .D(n8194), .CK(clk), .Q(reg_mem[477]) );
  DFF_X1 reg_mem_reg_196__4_ ( .D(n8193), .CK(clk), .Q(reg_mem[476]) );
  DFF_X1 reg_mem_reg_196__3_ ( .D(n8192), .CK(clk), .Q(reg_mem[475]) );
  DFF_X1 reg_mem_reg_196__2_ ( .D(n8191), .CK(clk), .Q(reg_mem[474]) );
  DFF_X1 reg_mem_reg_196__1_ ( .D(n8190), .CK(clk), .Q(reg_mem[473]) );
  DFF_X1 reg_mem_reg_196__0_ ( .D(n8189), .CK(clk), .Q(reg_mem[472]) );
  DFF_X1 reg_mem_reg_197__7_ ( .D(n7619), .CK(clk), .Q(reg_mem[471]) );
  DFF_X1 reg_mem_reg_197__6_ ( .D(n7618), .CK(clk), .Q(reg_mem[470]) );
  DFF_X1 reg_mem_reg_197__5_ ( .D(n7617), .CK(clk), .Q(reg_mem[469]) );
  DFF_X1 reg_mem_reg_197__4_ ( .D(n7616), .CK(clk), .Q(reg_mem[468]) );
  DFF_X1 reg_mem_reg_197__3_ ( .D(n7615), .CK(clk), .Q(reg_mem[467]) );
  DFF_X1 reg_mem_reg_197__2_ ( .D(n7614), .CK(clk), .Q(reg_mem[466]) );
  DFF_X1 reg_mem_reg_197__1_ ( .D(n7613), .CK(clk), .Q(reg_mem[465]) );
  DFF_X1 reg_mem_reg_197__0_ ( .D(n7612), .CK(clk), .Q(reg_mem[464]) );
  DFF_X1 reg_mem_reg_198__7_ ( .D(n8772), .CK(clk), .Q(reg_mem[463]) );
  DFF_X1 reg_mem_reg_198__6_ ( .D(n8771), .CK(clk), .Q(reg_mem[462]) );
  DFF_X1 reg_mem_reg_198__5_ ( .D(n8770), .CK(clk), .Q(reg_mem[461]) );
  DFF_X1 reg_mem_reg_198__4_ ( .D(n8769), .CK(clk), .Q(reg_mem[460]) );
  DFF_X1 reg_mem_reg_198__3_ ( .D(n8768), .CK(clk), .Q(reg_mem[459]) );
  DFF_X1 reg_mem_reg_198__2_ ( .D(n8767), .CK(clk), .Q(reg_mem[458]) );
  DFF_X1 reg_mem_reg_198__1_ ( .D(n8766), .CK(clk), .Q(reg_mem[457]) );
  DFF_X1 reg_mem_reg_198__0_ ( .D(n8765), .CK(clk), .Q(reg_mem[456]) );
  DFF_X1 reg_mem_reg_199__7_ ( .D(n7043), .CK(clk), .Q(reg_mem[455]) );
  DFF_X1 reg_mem_reg_199__6_ ( .D(n7042), .CK(clk), .Q(reg_mem[454]) );
  DFF_X1 reg_mem_reg_199__5_ ( .D(n7041), .CK(clk), .Q(reg_mem[453]) );
  DFF_X1 reg_mem_reg_199__4_ ( .D(n7040), .CK(clk), .Q(reg_mem[452]) );
  DFF_X1 reg_mem_reg_199__3_ ( .D(n7039), .CK(clk), .Q(reg_mem[451]) );
  DFF_X1 reg_mem_reg_199__2_ ( .D(n7038), .CK(clk), .Q(reg_mem[450]) );
  DFF_X1 reg_mem_reg_199__1_ ( .D(n7037), .CK(clk), .Q(reg_mem[449]) );
  DFF_X1 reg_mem_reg_199__0_ ( .D(n7036), .CK(clk), .Q(reg_mem[448]) );
  DFF_X1 reg_mem_reg_200__7_ ( .D(n8340), .CK(clk), .Q(reg_mem[447]) );
  DFF_X1 reg_mem_reg_200__6_ ( .D(n8339), .CK(clk), .Q(reg_mem[446]) );
  DFF_X1 reg_mem_reg_200__5_ ( .D(n8338), .CK(clk), .Q(reg_mem[445]) );
  DFF_X1 reg_mem_reg_200__4_ ( .D(n8337), .CK(clk), .Q(reg_mem[444]) );
  DFF_X1 reg_mem_reg_200__3_ ( .D(n8336), .CK(clk), .Q(reg_mem[443]) );
  DFF_X1 reg_mem_reg_200__2_ ( .D(n8335), .CK(clk), .Q(reg_mem[442]) );
  DFF_X1 reg_mem_reg_200__1_ ( .D(n8334), .CK(clk), .Q(reg_mem[441]) );
  DFF_X1 reg_mem_reg_200__0_ ( .D(n8333), .CK(clk), .Q(reg_mem[440]) );
  DFF_X1 reg_mem_reg_201__7_ ( .D(n7763), .CK(clk), .Q(reg_mem[439]) );
  DFF_X1 reg_mem_reg_201__6_ ( .D(n7762), .CK(clk), .Q(reg_mem[438]) );
  DFF_X1 reg_mem_reg_201__5_ ( .D(n7761), .CK(clk), .Q(reg_mem[437]) );
  DFF_X1 reg_mem_reg_201__4_ ( .D(n7760), .CK(clk), .Q(reg_mem[436]) );
  DFF_X1 reg_mem_reg_201__3_ ( .D(n7759), .CK(clk), .Q(reg_mem[435]) );
  DFF_X1 reg_mem_reg_201__2_ ( .D(n7758), .CK(clk), .Q(reg_mem[434]) );
  DFF_X1 reg_mem_reg_201__1_ ( .D(n7757), .CK(clk), .Q(reg_mem[433]) );
  DFF_X1 reg_mem_reg_201__0_ ( .D(n7756), .CK(clk), .Q(reg_mem[432]) );
  DFF_X1 reg_mem_reg_202__7_ ( .D(n8916), .CK(clk), .Q(reg_mem[431]) );
  DFF_X1 reg_mem_reg_202__6_ ( .D(n8915), .CK(clk), .Q(reg_mem[430]) );
  DFF_X1 reg_mem_reg_202__5_ ( .D(n8914), .CK(clk), .Q(reg_mem[429]) );
  DFF_X1 reg_mem_reg_202__4_ ( .D(n8913), .CK(clk), .Q(reg_mem[428]) );
  DFF_X1 reg_mem_reg_202__3_ ( .D(n8912), .CK(clk), .Q(reg_mem[427]) );
  DFF_X1 reg_mem_reg_202__2_ ( .D(n8911), .CK(clk), .Q(reg_mem[426]) );
  DFF_X1 reg_mem_reg_202__1_ ( .D(n8910), .CK(clk), .Q(reg_mem[425]) );
  DFF_X1 reg_mem_reg_202__0_ ( .D(n8909), .CK(clk), .Q(reg_mem[424]) );
  DFF_X1 reg_mem_reg_203__7_ ( .D(n7187), .CK(clk), .Q(reg_mem[423]) );
  DFF_X1 reg_mem_reg_203__6_ ( .D(n7186), .CK(clk), .Q(reg_mem[422]) );
  DFF_X1 reg_mem_reg_203__5_ ( .D(n7185), .CK(clk), .Q(reg_mem[421]) );
  DFF_X1 reg_mem_reg_203__4_ ( .D(n7184), .CK(clk), .Q(reg_mem[420]) );
  DFF_X1 reg_mem_reg_203__3_ ( .D(n7183), .CK(clk), .Q(reg_mem[419]) );
  DFF_X1 reg_mem_reg_203__2_ ( .D(n7182), .CK(clk), .Q(reg_mem[418]) );
  DFF_X1 reg_mem_reg_203__1_ ( .D(n7181), .CK(clk), .Q(reg_mem[417]) );
  DFF_X1 reg_mem_reg_203__0_ ( .D(n7180), .CK(clk), .Q(reg_mem[416]) );
  DFF_X1 reg_mem_reg_204__7_ ( .D(n8484), .CK(clk), .Q(reg_mem[415]) );
  DFF_X1 reg_mem_reg_204__6_ ( .D(n8483), .CK(clk), .Q(reg_mem[414]) );
  DFF_X1 reg_mem_reg_204__5_ ( .D(n8482), .CK(clk), .Q(reg_mem[413]) );
  DFF_X1 reg_mem_reg_204__4_ ( .D(n8481), .CK(clk), .Q(reg_mem[412]) );
  DFF_X1 reg_mem_reg_204__3_ ( .D(n8480), .CK(clk), .Q(reg_mem[411]) );
  DFF_X1 reg_mem_reg_204__2_ ( .D(n8479), .CK(clk), .Q(reg_mem[410]) );
  DFF_X1 reg_mem_reg_204__1_ ( .D(n8478), .CK(clk), .Q(reg_mem[409]) );
  DFF_X1 reg_mem_reg_204__0_ ( .D(n8477), .CK(clk), .Q(reg_mem[408]) );
  DFF_X1 reg_mem_reg_205__7_ ( .D(n7907), .CK(clk), .Q(reg_mem[407]) );
  DFF_X1 reg_mem_reg_205__6_ ( .D(n7906), .CK(clk), .Q(reg_mem[406]) );
  DFF_X1 reg_mem_reg_205__5_ ( .D(n7905), .CK(clk), .Q(reg_mem[405]) );
  DFF_X1 reg_mem_reg_205__4_ ( .D(n7904), .CK(clk), .Q(reg_mem[404]) );
  DFF_X1 reg_mem_reg_205__3_ ( .D(n7903), .CK(clk), .Q(reg_mem[403]) );
  DFF_X1 reg_mem_reg_205__2_ ( .D(n7902), .CK(clk), .Q(reg_mem[402]) );
  DFF_X1 reg_mem_reg_205__1_ ( .D(n7901), .CK(clk), .Q(reg_mem[401]) );
  DFF_X1 reg_mem_reg_205__0_ ( .D(n7900), .CK(clk), .Q(reg_mem[400]) );
  DFF_X1 reg_mem_reg_206__7_ ( .D(n9060), .CK(clk), .Q(reg_mem[399]) );
  DFF_X1 reg_mem_reg_206__6_ ( .D(n9059), .CK(clk), .Q(reg_mem[398]) );
  DFF_X1 reg_mem_reg_206__5_ ( .D(n9058), .CK(clk), .Q(reg_mem[397]) );
  DFF_X1 reg_mem_reg_206__4_ ( .D(n9057), .CK(clk), .Q(reg_mem[396]) );
  DFF_X1 reg_mem_reg_206__3_ ( .D(n9056), .CK(clk), .Q(reg_mem[395]) );
  DFF_X1 reg_mem_reg_206__2_ ( .D(n9055), .CK(clk), .Q(reg_mem[394]) );
  DFF_X1 reg_mem_reg_206__1_ ( .D(n9054), .CK(clk), .Q(reg_mem[393]) );
  DFF_X1 reg_mem_reg_206__0_ ( .D(n9053), .CK(clk), .Q(reg_mem[392]) );
  DFF_X1 reg_mem_reg_207__7_ ( .D(n7331), .CK(clk), .Q(reg_mem[391]) );
  DFF_X1 reg_mem_reg_207__6_ ( .D(n7330), .CK(clk), .Q(reg_mem[390]) );
  DFF_X1 reg_mem_reg_207__5_ ( .D(n7329), .CK(clk), .Q(reg_mem[389]) );
  DFF_X1 reg_mem_reg_207__4_ ( .D(n7328), .CK(clk), .Q(reg_mem[388]) );
  DFF_X1 reg_mem_reg_207__3_ ( .D(n7327), .CK(clk), .Q(reg_mem[387]) );
  DFF_X1 reg_mem_reg_207__2_ ( .D(n7326), .CK(clk), .Q(reg_mem[386]) );
  DFF_X1 reg_mem_reg_207__1_ ( .D(n7325), .CK(clk), .Q(reg_mem[385]) );
  DFF_X1 reg_mem_reg_207__0_ ( .D(n7324), .CK(clk), .Q(reg_mem[384]) );
  DFF_X1 reg_mem_reg_208__7_ ( .D(n8061), .CK(clk), .Q(reg_mem[383]) );
  DFF_X1 reg_mem_reg_208__6_ ( .D(n8060), .CK(clk), .Q(reg_mem[382]) );
  DFF_X1 reg_mem_reg_208__5_ ( .D(n8059), .CK(clk), .Q(reg_mem[381]) );
  DFF_X1 reg_mem_reg_208__4_ ( .D(n8058), .CK(clk), .Q(reg_mem[380]) );
  DFF_X1 reg_mem_reg_208__3_ ( .D(n8057), .CK(clk), .Q(reg_mem[379]) );
  DFF_X1 reg_mem_reg_208__2_ ( .D(n8056), .CK(clk), .Q(reg_mem[378]) );
  DFF_X1 reg_mem_reg_208__1_ ( .D(n8055), .CK(clk), .Q(reg_mem[377]) );
  DFF_X1 reg_mem_reg_208__0_ ( .D(n8054), .CK(clk), .Q(reg_mem[376]) );
  DFF_X1 reg_mem_reg_209__7_ ( .D(n7484), .CK(clk), .Q(reg_mem[375]) );
  DFF_X1 reg_mem_reg_209__6_ ( .D(n7483), .CK(clk), .Q(reg_mem[374]) );
  DFF_X1 reg_mem_reg_209__5_ ( .D(n7482), .CK(clk), .Q(reg_mem[373]) );
  DFF_X1 reg_mem_reg_209__4_ ( .D(n7481), .CK(clk), .Q(reg_mem[372]) );
  DFF_X1 reg_mem_reg_209__3_ ( .D(n7480), .CK(clk), .Q(reg_mem[371]) );
  DFF_X1 reg_mem_reg_209__2_ ( .D(n7479), .CK(clk), .Q(reg_mem[370]) );
  DFF_X1 reg_mem_reg_209__1_ ( .D(n7478), .CK(clk), .Q(reg_mem[369]) );
  DFF_X1 reg_mem_reg_209__0_ ( .D(n7477), .CK(clk), .Q(reg_mem[368]) );
  DFF_X1 reg_mem_reg_210__7_ ( .D(n8637), .CK(clk), .Q(reg_mem[367]) );
  DFF_X1 reg_mem_reg_210__6_ ( .D(n8636), .CK(clk), .Q(reg_mem[366]) );
  DFF_X1 reg_mem_reg_210__5_ ( .D(n8635), .CK(clk), .Q(reg_mem[365]) );
  DFF_X1 reg_mem_reg_210__4_ ( .D(n8634), .CK(clk), .Q(reg_mem[364]) );
  DFF_X1 reg_mem_reg_210__3_ ( .D(n8633), .CK(clk), .Q(reg_mem[363]) );
  DFF_X1 reg_mem_reg_210__2_ ( .D(n8632), .CK(clk), .Q(reg_mem[362]) );
  DFF_X1 reg_mem_reg_210__1_ ( .D(n8631), .CK(clk), .Q(reg_mem[361]) );
  DFF_X1 reg_mem_reg_210__0_ ( .D(n8630), .CK(clk), .Q(reg_mem[360]) );
  DFF_X1 reg_mem_reg_211__7_ ( .D(n6908), .CK(clk), .Q(reg_mem[359]) );
  DFF_X1 reg_mem_reg_211__6_ ( .D(n6907), .CK(clk), .Q(reg_mem[358]) );
  DFF_X1 reg_mem_reg_211__5_ ( .D(n6906), .CK(clk), .Q(reg_mem[357]) );
  DFF_X1 reg_mem_reg_211__4_ ( .D(n6905), .CK(clk), .Q(reg_mem[356]) );
  DFF_X1 reg_mem_reg_211__3_ ( .D(n6904), .CK(clk), .Q(reg_mem[355]) );
  DFF_X1 reg_mem_reg_211__2_ ( .D(n6903), .CK(clk), .Q(reg_mem[354]) );
  DFF_X1 reg_mem_reg_211__1_ ( .D(n6902), .CK(clk), .Q(reg_mem[353]) );
  DFF_X1 reg_mem_reg_211__0_ ( .D(n6901), .CK(clk), .Q(reg_mem[352]) );
  DFF_X1 reg_mem_reg_212__7_ ( .D(n8205), .CK(clk), .Q(reg_mem[351]) );
  DFF_X1 reg_mem_reg_212__6_ ( .D(n8204), .CK(clk), .Q(reg_mem[350]) );
  DFF_X1 reg_mem_reg_212__5_ ( .D(n8203), .CK(clk), .Q(reg_mem[349]) );
  DFF_X1 reg_mem_reg_212__4_ ( .D(n8202), .CK(clk), .Q(reg_mem[348]) );
  DFF_X1 reg_mem_reg_212__3_ ( .D(n8201), .CK(clk), .Q(reg_mem[347]) );
  DFF_X1 reg_mem_reg_212__2_ ( .D(n8200), .CK(clk), .Q(reg_mem[346]) );
  DFF_X1 reg_mem_reg_212__1_ ( .D(n8199), .CK(clk), .Q(reg_mem[345]) );
  DFF_X1 reg_mem_reg_212__0_ ( .D(n8198), .CK(clk), .Q(reg_mem[344]) );
  DFF_X1 reg_mem_reg_213__7_ ( .D(n7628), .CK(clk), .Q(reg_mem[343]) );
  DFF_X1 reg_mem_reg_213__6_ ( .D(n7627), .CK(clk), .Q(reg_mem[342]) );
  DFF_X1 reg_mem_reg_213__5_ ( .D(n7626), .CK(clk), .Q(reg_mem[341]) );
  DFF_X1 reg_mem_reg_213__4_ ( .D(n7625), .CK(clk), .Q(reg_mem[340]) );
  DFF_X1 reg_mem_reg_213__3_ ( .D(n7624), .CK(clk), .Q(reg_mem[339]) );
  DFF_X1 reg_mem_reg_213__2_ ( .D(n7623), .CK(clk), .Q(reg_mem[338]) );
  DFF_X1 reg_mem_reg_213__1_ ( .D(n7622), .CK(clk), .Q(reg_mem[337]) );
  DFF_X1 reg_mem_reg_213__0_ ( .D(n7621), .CK(clk), .Q(reg_mem[336]) );
  DFF_X1 reg_mem_reg_214__7_ ( .D(n8781), .CK(clk), .Q(reg_mem[335]) );
  DFF_X1 reg_mem_reg_214__6_ ( .D(n8780), .CK(clk), .Q(reg_mem[334]) );
  DFF_X1 reg_mem_reg_214__5_ ( .D(n8779), .CK(clk), .Q(reg_mem[333]) );
  DFF_X1 reg_mem_reg_214__4_ ( .D(n8778), .CK(clk), .Q(reg_mem[332]) );
  DFF_X1 reg_mem_reg_214__3_ ( .D(n8777), .CK(clk), .Q(reg_mem[331]) );
  DFF_X1 reg_mem_reg_214__2_ ( .D(n8776), .CK(clk), .Q(reg_mem[330]) );
  DFF_X1 reg_mem_reg_214__1_ ( .D(n8775), .CK(clk), .Q(reg_mem[329]) );
  DFF_X1 reg_mem_reg_214__0_ ( .D(n8774), .CK(clk), .Q(reg_mem[328]) );
  DFF_X1 reg_mem_reg_215__7_ ( .D(n7052), .CK(clk), .Q(reg_mem[327]) );
  DFF_X1 reg_mem_reg_215__6_ ( .D(n7051), .CK(clk), .Q(reg_mem[326]) );
  DFF_X1 reg_mem_reg_215__5_ ( .D(n7050), .CK(clk), .Q(reg_mem[325]) );
  DFF_X1 reg_mem_reg_215__4_ ( .D(n7049), .CK(clk), .Q(reg_mem[324]) );
  DFF_X1 reg_mem_reg_215__3_ ( .D(n7048), .CK(clk), .Q(reg_mem[323]) );
  DFF_X1 reg_mem_reg_215__2_ ( .D(n7047), .CK(clk), .Q(reg_mem[322]) );
  DFF_X1 reg_mem_reg_215__1_ ( .D(n7046), .CK(clk), .Q(reg_mem[321]) );
  DFF_X1 reg_mem_reg_215__0_ ( .D(n7045), .CK(clk), .Q(reg_mem[320]) );
  DFF_X1 reg_mem_reg_216__7_ ( .D(n8349), .CK(clk), .Q(reg_mem[319]) );
  DFF_X1 reg_mem_reg_216__6_ ( .D(n8348), .CK(clk), .Q(reg_mem[318]) );
  DFF_X1 reg_mem_reg_216__5_ ( .D(n8347), .CK(clk), .Q(reg_mem[317]) );
  DFF_X1 reg_mem_reg_216__4_ ( .D(n8346), .CK(clk), .Q(reg_mem[316]) );
  DFF_X1 reg_mem_reg_216__3_ ( .D(n8345), .CK(clk), .Q(reg_mem[315]) );
  DFF_X1 reg_mem_reg_216__2_ ( .D(n8344), .CK(clk), .Q(reg_mem[314]) );
  DFF_X1 reg_mem_reg_216__1_ ( .D(n8343), .CK(clk), .Q(reg_mem[313]) );
  DFF_X1 reg_mem_reg_216__0_ ( .D(n8342), .CK(clk), .Q(reg_mem[312]) );
  DFF_X1 reg_mem_reg_217__7_ ( .D(n7772), .CK(clk), .Q(reg_mem[311]) );
  DFF_X1 reg_mem_reg_217__6_ ( .D(n7771), .CK(clk), .Q(reg_mem[310]) );
  DFF_X1 reg_mem_reg_217__5_ ( .D(n7770), .CK(clk), .Q(reg_mem[309]) );
  DFF_X1 reg_mem_reg_217__4_ ( .D(n7769), .CK(clk), .Q(reg_mem[308]) );
  DFF_X1 reg_mem_reg_217__3_ ( .D(n7768), .CK(clk), .Q(reg_mem[307]) );
  DFF_X1 reg_mem_reg_217__2_ ( .D(n7767), .CK(clk), .Q(reg_mem[306]) );
  DFF_X1 reg_mem_reg_217__1_ ( .D(n7766), .CK(clk), .Q(reg_mem[305]) );
  DFF_X1 reg_mem_reg_217__0_ ( .D(n7765), .CK(clk), .Q(reg_mem[304]) );
  DFF_X1 reg_mem_reg_218__7_ ( .D(n8925), .CK(clk), .Q(reg_mem[303]) );
  DFF_X1 reg_mem_reg_218__6_ ( .D(n8924), .CK(clk), .Q(reg_mem[302]) );
  DFF_X1 reg_mem_reg_218__5_ ( .D(n8923), .CK(clk), .Q(reg_mem[301]) );
  DFF_X1 reg_mem_reg_218__4_ ( .D(n8922), .CK(clk), .Q(reg_mem[300]) );
  DFF_X1 reg_mem_reg_218__3_ ( .D(n8921), .CK(clk), .Q(reg_mem[299]) );
  DFF_X1 reg_mem_reg_218__2_ ( .D(n8920), .CK(clk), .Q(reg_mem[298]) );
  DFF_X1 reg_mem_reg_218__1_ ( .D(n8919), .CK(clk), .Q(reg_mem[297]) );
  DFF_X1 reg_mem_reg_218__0_ ( .D(n8918), .CK(clk), .Q(reg_mem[296]) );
  DFF_X1 reg_mem_reg_219__7_ ( .D(n7196), .CK(clk), .Q(reg_mem[295]) );
  DFF_X1 reg_mem_reg_219__6_ ( .D(n7195), .CK(clk), .Q(reg_mem[294]) );
  DFF_X1 reg_mem_reg_219__5_ ( .D(n7194), .CK(clk), .Q(reg_mem[293]) );
  DFF_X1 reg_mem_reg_219__4_ ( .D(n7193), .CK(clk), .Q(reg_mem[292]) );
  DFF_X1 reg_mem_reg_219__3_ ( .D(n7192), .CK(clk), .Q(reg_mem[291]) );
  DFF_X1 reg_mem_reg_219__2_ ( .D(n7191), .CK(clk), .Q(reg_mem[290]) );
  DFF_X1 reg_mem_reg_219__1_ ( .D(n7190), .CK(clk), .Q(reg_mem[289]) );
  DFF_X1 reg_mem_reg_219__0_ ( .D(n7189), .CK(clk), .Q(reg_mem[288]) );
  DFF_X1 reg_mem_reg_220__7_ ( .D(n8493), .CK(clk), .Q(reg_mem[287]) );
  DFF_X1 reg_mem_reg_220__6_ ( .D(n8492), .CK(clk), .Q(reg_mem[286]) );
  DFF_X1 reg_mem_reg_220__5_ ( .D(n8491), .CK(clk), .Q(reg_mem[285]) );
  DFF_X1 reg_mem_reg_220__4_ ( .D(n8490), .CK(clk), .Q(reg_mem[284]) );
  DFF_X1 reg_mem_reg_220__3_ ( .D(n8489), .CK(clk), .Q(reg_mem[283]) );
  DFF_X1 reg_mem_reg_220__2_ ( .D(n8488), .CK(clk), .Q(reg_mem[282]) );
  DFF_X1 reg_mem_reg_220__1_ ( .D(n8487), .CK(clk), .Q(reg_mem[281]) );
  DFF_X1 reg_mem_reg_220__0_ ( .D(n8486), .CK(clk), .Q(reg_mem[280]) );
  DFF_X1 reg_mem_reg_221__7_ ( .D(n7916), .CK(clk), .Q(reg_mem[279]) );
  DFF_X1 reg_mem_reg_221__6_ ( .D(n7915), .CK(clk), .Q(reg_mem[278]) );
  DFF_X1 reg_mem_reg_221__5_ ( .D(n7914), .CK(clk), .Q(reg_mem[277]) );
  DFF_X1 reg_mem_reg_221__4_ ( .D(n7913), .CK(clk), .Q(reg_mem[276]) );
  DFF_X1 reg_mem_reg_221__3_ ( .D(n7912), .CK(clk), .Q(reg_mem[275]) );
  DFF_X1 reg_mem_reg_221__2_ ( .D(n7911), .CK(clk), .Q(reg_mem[274]) );
  DFF_X1 reg_mem_reg_221__1_ ( .D(n7910), .CK(clk), .Q(reg_mem[273]) );
  DFF_X1 reg_mem_reg_221__0_ ( .D(n7909), .CK(clk), .Q(reg_mem[272]) );
  DFF_X1 reg_mem_reg_222__7_ ( .D(n9069), .CK(clk), .Q(reg_mem[271]) );
  DFF_X1 reg_mem_reg_222__6_ ( .D(n9068), .CK(clk), .Q(reg_mem[270]) );
  DFF_X1 reg_mem_reg_222__5_ ( .D(n9067), .CK(clk), .Q(reg_mem[269]) );
  DFF_X1 reg_mem_reg_222__4_ ( .D(n9066), .CK(clk), .Q(reg_mem[268]) );
  DFF_X1 reg_mem_reg_222__3_ ( .D(n9065), .CK(clk), .Q(reg_mem[267]) );
  DFF_X1 reg_mem_reg_222__2_ ( .D(n9064), .CK(clk), .Q(reg_mem[266]) );
  DFF_X1 reg_mem_reg_222__1_ ( .D(n9063), .CK(clk), .Q(reg_mem[265]) );
  DFF_X1 reg_mem_reg_222__0_ ( .D(n9062), .CK(clk), .Q(reg_mem[264]) );
  DFF_X1 reg_mem_reg_223__7_ ( .D(n7340), .CK(clk), .Q(reg_mem[263]) );
  DFF_X1 reg_mem_reg_223__6_ ( .D(n7339), .CK(clk), .Q(reg_mem[262]) );
  DFF_X1 reg_mem_reg_223__5_ ( .D(n7338), .CK(clk), .Q(reg_mem[261]) );
  DFF_X1 reg_mem_reg_223__4_ ( .D(n7337), .CK(clk), .Q(reg_mem[260]) );
  DFF_X1 reg_mem_reg_223__3_ ( .D(n7336), .CK(clk), .Q(reg_mem[259]) );
  DFF_X1 reg_mem_reg_223__2_ ( .D(n7335), .CK(clk), .Q(reg_mem[258]) );
  DFF_X1 reg_mem_reg_223__1_ ( .D(n7334), .CK(clk), .Q(reg_mem[257]) );
  DFF_X1 reg_mem_reg_223__0_ ( .D(n7333), .CK(clk), .Q(reg_mem[256]) );
  DFF_X1 reg_mem_reg_224__7_ ( .D(n8070), .CK(clk), .Q(reg_mem[255]) );
  DFF_X1 reg_mem_reg_224__6_ ( .D(n8069), .CK(clk), .Q(reg_mem[254]) );
  DFF_X1 reg_mem_reg_224__5_ ( .D(n8068), .CK(clk), .Q(reg_mem[253]) );
  DFF_X1 reg_mem_reg_224__4_ ( .D(n8067), .CK(clk), .Q(reg_mem[252]) );
  DFF_X1 reg_mem_reg_224__3_ ( .D(n8066), .CK(clk), .Q(reg_mem[251]) );
  DFF_X1 reg_mem_reg_224__2_ ( .D(n8065), .CK(clk), .Q(reg_mem[250]) );
  DFF_X1 reg_mem_reg_224__1_ ( .D(n8064), .CK(clk), .Q(reg_mem[249]) );
  DFF_X1 reg_mem_reg_224__0_ ( .D(n8063), .CK(clk), .Q(reg_mem[248]) );
  DFF_X1 reg_mem_reg_225__7_ ( .D(n7493), .CK(clk), .Q(reg_mem[247]) );
  DFF_X1 reg_mem_reg_225__6_ ( .D(n7492), .CK(clk), .Q(reg_mem[246]) );
  DFF_X1 reg_mem_reg_225__5_ ( .D(n7491), .CK(clk), .Q(reg_mem[245]) );
  DFF_X1 reg_mem_reg_225__4_ ( .D(n7490), .CK(clk), .Q(reg_mem[244]) );
  DFF_X1 reg_mem_reg_225__3_ ( .D(n7489), .CK(clk), .Q(reg_mem[243]) );
  DFF_X1 reg_mem_reg_225__2_ ( .D(n7488), .CK(clk), .Q(reg_mem[242]) );
  DFF_X1 reg_mem_reg_225__1_ ( .D(n7487), .CK(clk), .Q(reg_mem[241]) );
  DFF_X1 reg_mem_reg_225__0_ ( .D(n7486), .CK(clk), .Q(reg_mem[240]) );
  DFF_X1 reg_mem_reg_226__7_ ( .D(n8646), .CK(clk), .Q(reg_mem[239]) );
  DFF_X1 reg_mem_reg_226__6_ ( .D(n8645), .CK(clk), .Q(reg_mem[238]) );
  DFF_X1 reg_mem_reg_226__5_ ( .D(n8644), .CK(clk), .Q(reg_mem[237]) );
  DFF_X1 reg_mem_reg_226__4_ ( .D(n8643), .CK(clk), .Q(reg_mem[236]) );
  DFF_X1 reg_mem_reg_226__3_ ( .D(n8642), .CK(clk), .Q(reg_mem[235]) );
  DFF_X1 reg_mem_reg_226__2_ ( .D(n8641), .CK(clk), .Q(reg_mem[234]) );
  DFF_X1 reg_mem_reg_226__1_ ( .D(n8640), .CK(clk), .Q(reg_mem[233]) );
  DFF_X1 reg_mem_reg_226__0_ ( .D(n8639), .CK(clk), .Q(reg_mem[232]) );
  DFF_X1 reg_mem_reg_227__7_ ( .D(n6917), .CK(clk), .Q(reg_mem[231]) );
  DFF_X1 reg_mem_reg_227__6_ ( .D(n6916), .CK(clk), .Q(reg_mem[230]) );
  DFF_X1 reg_mem_reg_227__5_ ( .D(n6915), .CK(clk), .Q(reg_mem[229]) );
  DFF_X1 reg_mem_reg_227__4_ ( .D(n6914), .CK(clk), .Q(reg_mem[228]) );
  DFF_X1 reg_mem_reg_227__3_ ( .D(n6913), .CK(clk), .Q(reg_mem[227]) );
  DFF_X1 reg_mem_reg_227__2_ ( .D(n6912), .CK(clk), .Q(reg_mem[226]) );
  DFF_X1 reg_mem_reg_227__1_ ( .D(n6911), .CK(clk), .Q(reg_mem[225]) );
  DFF_X1 reg_mem_reg_227__0_ ( .D(n6910), .CK(clk), .Q(reg_mem[224]) );
  DFF_X1 reg_mem_reg_228__7_ ( .D(n8214), .CK(clk), .Q(reg_mem[223]) );
  DFF_X1 reg_mem_reg_228__6_ ( .D(n8213), .CK(clk), .Q(reg_mem[222]) );
  DFF_X1 reg_mem_reg_228__5_ ( .D(n8212), .CK(clk), .Q(reg_mem[221]) );
  DFF_X1 reg_mem_reg_228__4_ ( .D(n8211), .CK(clk), .Q(reg_mem[220]) );
  DFF_X1 reg_mem_reg_228__3_ ( .D(n8210), .CK(clk), .Q(reg_mem[219]) );
  DFF_X1 reg_mem_reg_228__2_ ( .D(n8209), .CK(clk), .Q(reg_mem[218]) );
  DFF_X1 reg_mem_reg_228__1_ ( .D(n8208), .CK(clk), .Q(reg_mem[217]) );
  DFF_X1 reg_mem_reg_228__0_ ( .D(n8207), .CK(clk), .Q(reg_mem[216]) );
  DFF_X1 reg_mem_reg_229__7_ ( .D(n7637), .CK(clk), .Q(reg_mem[215]) );
  DFF_X1 reg_mem_reg_229__6_ ( .D(n7636), .CK(clk), .Q(reg_mem[214]) );
  DFF_X1 reg_mem_reg_229__5_ ( .D(n7635), .CK(clk), .Q(reg_mem[213]) );
  DFF_X1 reg_mem_reg_229__4_ ( .D(n7634), .CK(clk), .Q(reg_mem[212]) );
  DFF_X1 reg_mem_reg_229__3_ ( .D(n7633), .CK(clk), .Q(reg_mem[211]) );
  DFF_X1 reg_mem_reg_229__2_ ( .D(n7632), .CK(clk), .Q(reg_mem[210]) );
  DFF_X1 reg_mem_reg_229__1_ ( .D(n7631), .CK(clk), .Q(reg_mem[209]) );
  DFF_X1 reg_mem_reg_229__0_ ( .D(n7630), .CK(clk), .Q(reg_mem[208]) );
  DFF_X1 reg_mem_reg_230__7_ ( .D(n8790), .CK(clk), .Q(reg_mem[207]) );
  DFF_X1 reg_mem_reg_230__6_ ( .D(n8789), .CK(clk), .Q(reg_mem[206]) );
  DFF_X1 reg_mem_reg_230__5_ ( .D(n8788), .CK(clk), .Q(reg_mem[205]) );
  DFF_X1 reg_mem_reg_230__4_ ( .D(n8787), .CK(clk), .Q(reg_mem[204]) );
  DFF_X1 reg_mem_reg_230__3_ ( .D(n8786), .CK(clk), .Q(reg_mem[203]) );
  DFF_X1 reg_mem_reg_230__2_ ( .D(n8785), .CK(clk), .Q(reg_mem[202]) );
  DFF_X1 reg_mem_reg_230__1_ ( .D(n8784), .CK(clk), .Q(reg_mem[201]) );
  DFF_X1 reg_mem_reg_230__0_ ( .D(n8783), .CK(clk), .Q(reg_mem[200]) );
  DFF_X1 reg_mem_reg_231__7_ ( .D(n7061), .CK(clk), .Q(reg_mem[199]) );
  DFF_X1 reg_mem_reg_231__6_ ( .D(n7060), .CK(clk), .Q(reg_mem[198]) );
  DFF_X1 reg_mem_reg_231__5_ ( .D(n7059), .CK(clk), .Q(reg_mem[197]) );
  DFF_X1 reg_mem_reg_231__4_ ( .D(n7058), .CK(clk), .Q(reg_mem[196]) );
  DFF_X1 reg_mem_reg_231__3_ ( .D(n7057), .CK(clk), .Q(reg_mem[195]) );
  DFF_X1 reg_mem_reg_231__2_ ( .D(n7056), .CK(clk), .Q(reg_mem[194]) );
  DFF_X1 reg_mem_reg_231__1_ ( .D(n7055), .CK(clk), .Q(reg_mem[193]) );
  DFF_X1 reg_mem_reg_231__0_ ( .D(n7054), .CK(clk), .Q(reg_mem[192]) );
  DFF_X1 reg_mem_reg_232__7_ ( .D(n8358), .CK(clk), .Q(reg_mem[191]) );
  DFF_X1 reg_mem_reg_232__6_ ( .D(n8357), .CK(clk), .Q(reg_mem[190]) );
  DFF_X1 reg_mem_reg_232__5_ ( .D(n8356), .CK(clk), .Q(reg_mem[189]) );
  DFF_X1 reg_mem_reg_232__4_ ( .D(n8355), .CK(clk), .Q(reg_mem[188]) );
  DFF_X1 reg_mem_reg_232__3_ ( .D(n8354), .CK(clk), .Q(reg_mem[187]) );
  DFF_X1 reg_mem_reg_232__2_ ( .D(n8353), .CK(clk), .Q(reg_mem[186]) );
  DFF_X1 reg_mem_reg_232__1_ ( .D(n8352), .CK(clk), .Q(reg_mem[185]) );
  DFF_X1 reg_mem_reg_232__0_ ( .D(n8351), .CK(clk), .Q(reg_mem[184]) );
  DFF_X1 reg_mem_reg_233__7_ ( .D(n7781), .CK(clk), .Q(reg_mem[183]) );
  DFF_X1 reg_mem_reg_233__6_ ( .D(n7780), .CK(clk), .Q(reg_mem[182]) );
  DFF_X1 reg_mem_reg_233__5_ ( .D(n7779), .CK(clk), .Q(reg_mem[181]) );
  DFF_X1 reg_mem_reg_233__4_ ( .D(n7778), .CK(clk), .Q(reg_mem[180]) );
  DFF_X1 reg_mem_reg_233__3_ ( .D(n7777), .CK(clk), .Q(reg_mem[179]) );
  DFF_X1 reg_mem_reg_233__2_ ( .D(n7776), .CK(clk), .Q(reg_mem[178]) );
  DFF_X1 reg_mem_reg_233__1_ ( .D(n7775), .CK(clk), .Q(reg_mem[177]) );
  DFF_X1 reg_mem_reg_233__0_ ( .D(n7774), .CK(clk), .Q(reg_mem[176]) );
  DFF_X1 reg_mem_reg_234__7_ ( .D(n8934), .CK(clk), .Q(reg_mem[175]) );
  DFF_X1 reg_mem_reg_234__6_ ( .D(n8933), .CK(clk), .Q(reg_mem[174]) );
  DFF_X1 reg_mem_reg_234__5_ ( .D(n8932), .CK(clk), .Q(reg_mem[173]) );
  DFF_X1 reg_mem_reg_234__4_ ( .D(n8931), .CK(clk), .Q(reg_mem[172]) );
  DFF_X1 reg_mem_reg_234__3_ ( .D(n8930), .CK(clk), .Q(reg_mem[171]) );
  DFF_X1 reg_mem_reg_234__2_ ( .D(n8929), .CK(clk), .Q(reg_mem[170]) );
  DFF_X1 reg_mem_reg_234__1_ ( .D(n8928), .CK(clk), .Q(reg_mem[169]) );
  DFF_X1 reg_mem_reg_234__0_ ( .D(n8927), .CK(clk), .Q(reg_mem[168]) );
  DFF_X1 reg_mem_reg_235__7_ ( .D(n7205), .CK(clk), .Q(reg_mem[167]) );
  DFF_X1 reg_mem_reg_235__6_ ( .D(n7204), .CK(clk), .Q(reg_mem[166]) );
  DFF_X1 reg_mem_reg_235__5_ ( .D(n7203), .CK(clk), .Q(reg_mem[165]) );
  DFF_X1 reg_mem_reg_235__4_ ( .D(n7202), .CK(clk), .Q(reg_mem[164]) );
  DFF_X1 reg_mem_reg_235__3_ ( .D(n7201), .CK(clk), .Q(reg_mem[163]) );
  DFF_X1 reg_mem_reg_235__2_ ( .D(n7200), .CK(clk), .Q(reg_mem[162]) );
  DFF_X1 reg_mem_reg_235__1_ ( .D(n7199), .CK(clk), .Q(reg_mem[161]) );
  DFF_X1 reg_mem_reg_235__0_ ( .D(n7198), .CK(clk), .Q(reg_mem[160]) );
  DFF_X1 reg_mem_reg_236__7_ ( .D(n8502), .CK(clk), .Q(reg_mem[159]) );
  DFF_X1 reg_mem_reg_236__6_ ( .D(n8501), .CK(clk), .Q(reg_mem[158]) );
  DFF_X1 reg_mem_reg_236__5_ ( .D(n8500), .CK(clk), .Q(reg_mem[157]) );
  DFF_X1 reg_mem_reg_236__4_ ( .D(n8499), .CK(clk), .Q(reg_mem[156]) );
  DFF_X1 reg_mem_reg_236__3_ ( .D(n8498), .CK(clk), .Q(reg_mem[155]) );
  DFF_X1 reg_mem_reg_236__2_ ( .D(n8497), .CK(clk), .Q(reg_mem[154]) );
  DFF_X1 reg_mem_reg_236__1_ ( .D(n8496), .CK(clk), .Q(reg_mem[153]) );
  DFF_X1 reg_mem_reg_236__0_ ( .D(n8495), .CK(clk), .Q(reg_mem[152]) );
  DFF_X1 reg_mem_reg_237__7_ ( .D(n7925), .CK(clk), .Q(reg_mem[151]) );
  DFF_X1 reg_mem_reg_237__6_ ( .D(n7924), .CK(clk), .Q(reg_mem[150]) );
  DFF_X1 reg_mem_reg_237__5_ ( .D(n7923), .CK(clk), .Q(reg_mem[149]) );
  DFF_X1 reg_mem_reg_237__4_ ( .D(n7922), .CK(clk), .Q(reg_mem[148]) );
  DFF_X1 reg_mem_reg_237__3_ ( .D(n7921), .CK(clk), .Q(reg_mem[147]) );
  DFF_X1 reg_mem_reg_237__2_ ( .D(n7920), .CK(clk), .Q(reg_mem[146]) );
  DFF_X1 reg_mem_reg_237__1_ ( .D(n7919), .CK(clk), .Q(reg_mem[145]) );
  DFF_X1 reg_mem_reg_237__0_ ( .D(n7918), .CK(clk), .Q(reg_mem[144]) );
  DFF_X1 reg_mem_reg_238__7_ ( .D(n9078), .CK(clk), .Q(reg_mem[143]) );
  DFF_X1 reg_mem_reg_238__6_ ( .D(n9077), .CK(clk), .Q(reg_mem[142]) );
  DFF_X1 reg_mem_reg_238__5_ ( .D(n9076), .CK(clk), .Q(reg_mem[141]) );
  DFF_X1 reg_mem_reg_238__4_ ( .D(n9075), .CK(clk), .Q(reg_mem[140]) );
  DFF_X1 reg_mem_reg_238__3_ ( .D(n9074), .CK(clk), .Q(reg_mem[139]) );
  DFF_X1 reg_mem_reg_238__2_ ( .D(n9073), .CK(clk), .Q(reg_mem[138]) );
  DFF_X1 reg_mem_reg_238__1_ ( .D(n9072), .CK(clk), .Q(reg_mem[137]) );
  DFF_X1 reg_mem_reg_238__0_ ( .D(n9071), .CK(clk), .Q(reg_mem[136]) );
  DFF_X1 reg_mem_reg_239__7_ ( .D(n7349), .CK(clk), .Q(reg_mem[135]) );
  DFF_X1 reg_mem_reg_239__6_ ( .D(n7348), .CK(clk), .Q(reg_mem[134]) );
  DFF_X1 reg_mem_reg_239__5_ ( .D(n7347), .CK(clk), .Q(reg_mem[133]) );
  DFF_X1 reg_mem_reg_239__4_ ( .D(n7346), .CK(clk), .Q(reg_mem[132]) );
  DFF_X1 reg_mem_reg_239__3_ ( .D(n7345), .CK(clk), .Q(reg_mem[131]) );
  DFF_X1 reg_mem_reg_239__2_ ( .D(n7344), .CK(clk), .Q(reg_mem[130]) );
  DFF_X1 reg_mem_reg_239__1_ ( .D(n7343), .CK(clk), .Q(reg_mem[129]) );
  DFF_X1 reg_mem_reg_239__0_ ( .D(n7342), .CK(clk), .Q(reg_mem[128]) );
  DFF_X1 reg_mem_reg_240__7_ ( .D(n8079), .CK(clk), .Q(reg_mem[127]) );
  DFF_X1 reg_mem_reg_240__6_ ( .D(n8078), .CK(clk), .Q(reg_mem[126]) );
  DFF_X1 reg_mem_reg_240__5_ ( .D(n8077), .CK(clk), .Q(reg_mem[125]) );
  DFF_X1 reg_mem_reg_240__4_ ( .D(n8076), .CK(clk), .Q(reg_mem[124]) );
  DFF_X1 reg_mem_reg_240__3_ ( .D(n8075), .CK(clk), .Q(reg_mem[123]) );
  DFF_X1 reg_mem_reg_240__2_ ( .D(n8074), .CK(clk), .Q(reg_mem[122]) );
  DFF_X1 reg_mem_reg_240__1_ ( .D(n8073), .CK(clk), .Q(reg_mem[121]) );
  DFF_X1 reg_mem_reg_240__0_ ( .D(n8072), .CK(clk), .Q(reg_mem[120]) );
  DFF_X1 reg_mem_reg_241__7_ ( .D(n7502), .CK(clk), .Q(reg_mem[119]) );
  DFF_X1 reg_mem_reg_241__6_ ( .D(n7501), .CK(clk), .Q(reg_mem[118]) );
  DFF_X1 reg_mem_reg_241__5_ ( .D(n7500), .CK(clk), .Q(reg_mem[117]) );
  DFF_X1 reg_mem_reg_241__4_ ( .D(n7499), .CK(clk), .Q(reg_mem[116]) );
  DFF_X1 reg_mem_reg_241__3_ ( .D(n7498), .CK(clk), .Q(reg_mem[115]) );
  DFF_X1 reg_mem_reg_241__2_ ( .D(n7497), .CK(clk), .Q(reg_mem[114]) );
  DFF_X1 reg_mem_reg_241__1_ ( .D(n7496), .CK(clk), .Q(reg_mem[113]) );
  DFF_X1 reg_mem_reg_241__0_ ( .D(n7495), .CK(clk), .Q(reg_mem[112]) );
  DFF_X1 reg_mem_reg_242__7_ ( .D(n8655), .CK(clk), .Q(reg_mem[111]) );
  DFF_X1 reg_mem_reg_242__6_ ( .D(n8654), .CK(clk), .Q(reg_mem[110]) );
  DFF_X1 reg_mem_reg_242__5_ ( .D(n8653), .CK(clk), .Q(reg_mem[109]) );
  DFF_X1 reg_mem_reg_242__4_ ( .D(n8652), .CK(clk), .Q(reg_mem[108]) );
  DFF_X1 reg_mem_reg_242__3_ ( .D(n8651), .CK(clk), .Q(reg_mem[107]) );
  DFF_X1 reg_mem_reg_242__2_ ( .D(n8650), .CK(clk), .Q(reg_mem[106]) );
  DFF_X1 reg_mem_reg_242__1_ ( .D(n8649), .CK(clk), .Q(reg_mem[105]) );
  DFF_X1 reg_mem_reg_242__0_ ( .D(n8648), .CK(clk), .Q(reg_mem[104]) );
  DFF_X1 reg_mem_reg_243__7_ ( .D(n6926), .CK(clk), .Q(reg_mem[103]) );
  DFF_X1 reg_mem_reg_243__6_ ( .D(n6925), .CK(clk), .Q(reg_mem[102]) );
  DFF_X1 reg_mem_reg_243__5_ ( .D(n6924), .CK(clk), .Q(reg_mem[101]) );
  DFF_X1 reg_mem_reg_243__4_ ( .D(n6923), .CK(clk), .Q(reg_mem[100]) );
  DFF_X1 reg_mem_reg_243__3_ ( .D(n6922), .CK(clk), .Q(reg_mem[99]) );
  DFF_X1 reg_mem_reg_243__2_ ( .D(n6921), .CK(clk), .Q(reg_mem[98]) );
  DFF_X1 reg_mem_reg_243__1_ ( .D(n6920), .CK(clk), .Q(reg_mem[97]) );
  DFF_X1 reg_mem_reg_243__0_ ( .D(n6919), .CK(clk), .Q(reg_mem[96]) );
  DFF_X1 reg_mem_reg_244__7_ ( .D(n8223), .CK(clk), .Q(reg_mem[95]) );
  DFF_X1 reg_mem_reg_244__6_ ( .D(n8222), .CK(clk), .Q(reg_mem[94]) );
  DFF_X1 reg_mem_reg_244__5_ ( .D(n8221), .CK(clk), .Q(reg_mem[93]) );
  DFF_X1 reg_mem_reg_244__4_ ( .D(n8220), .CK(clk), .Q(reg_mem[92]) );
  DFF_X1 reg_mem_reg_244__3_ ( .D(n8219), .CK(clk), .Q(reg_mem[91]) );
  DFF_X1 reg_mem_reg_244__2_ ( .D(n8218), .CK(clk), .Q(reg_mem[90]) );
  DFF_X1 reg_mem_reg_244__1_ ( .D(n8217), .CK(clk), .Q(reg_mem[89]) );
  DFF_X1 reg_mem_reg_244__0_ ( .D(n8216), .CK(clk), .Q(reg_mem[88]) );
  DFF_X1 reg_mem_reg_245__7_ ( .D(n7646), .CK(clk), .Q(reg_mem[87]) );
  DFF_X1 reg_mem_reg_245__6_ ( .D(n7645), .CK(clk), .Q(reg_mem[86]) );
  DFF_X1 reg_mem_reg_245__5_ ( .D(n7644), .CK(clk), .Q(reg_mem[85]) );
  DFF_X1 reg_mem_reg_245__4_ ( .D(n7643), .CK(clk), .Q(reg_mem[84]) );
  DFF_X1 reg_mem_reg_245__3_ ( .D(n7642), .CK(clk), .Q(reg_mem[83]) );
  DFF_X1 reg_mem_reg_245__2_ ( .D(n7641), .CK(clk), .Q(reg_mem[82]) );
  DFF_X1 reg_mem_reg_245__1_ ( .D(n7640), .CK(clk), .Q(reg_mem[81]) );
  DFF_X1 reg_mem_reg_245__0_ ( .D(n7639), .CK(clk), .Q(reg_mem[80]) );
  DFF_X1 reg_mem_reg_246__7_ ( .D(n8799), .CK(clk), .Q(reg_mem[79]) );
  DFF_X1 reg_mem_reg_246__6_ ( .D(n8798), .CK(clk), .Q(reg_mem[78]) );
  DFF_X1 reg_mem_reg_246__5_ ( .D(n8797), .CK(clk), .Q(reg_mem[77]) );
  DFF_X1 reg_mem_reg_246__4_ ( .D(n8796), .CK(clk), .Q(reg_mem[76]) );
  DFF_X1 reg_mem_reg_246__3_ ( .D(n8795), .CK(clk), .Q(reg_mem[75]) );
  DFF_X1 reg_mem_reg_246__2_ ( .D(n8794), .CK(clk), .Q(reg_mem[74]) );
  DFF_X1 reg_mem_reg_246__1_ ( .D(n8793), .CK(clk), .Q(reg_mem[73]) );
  DFF_X1 reg_mem_reg_246__0_ ( .D(n8792), .CK(clk), .Q(reg_mem[72]) );
  DFF_X1 reg_mem_reg_247__7_ ( .D(n7070), .CK(clk), .Q(reg_mem[71]) );
  DFF_X1 reg_mem_reg_247__6_ ( .D(n7069), .CK(clk), .Q(reg_mem[70]) );
  DFF_X1 reg_mem_reg_247__5_ ( .D(n7068), .CK(clk), .Q(reg_mem[69]) );
  DFF_X1 reg_mem_reg_247__4_ ( .D(n7067), .CK(clk), .Q(reg_mem[68]) );
  DFF_X1 reg_mem_reg_247__3_ ( .D(n7066), .CK(clk), .Q(reg_mem[67]) );
  DFF_X1 reg_mem_reg_247__2_ ( .D(n7065), .CK(clk), .Q(reg_mem[66]) );
  DFF_X1 reg_mem_reg_247__1_ ( .D(n7064), .CK(clk), .Q(reg_mem[65]) );
  DFF_X1 reg_mem_reg_247__0_ ( .D(n7063), .CK(clk), .Q(reg_mem[64]) );
  DFF_X1 reg_mem_reg_248__7_ ( .D(n8367), .CK(clk), .Q(reg_mem[63]) );
  DFF_X1 reg_mem_reg_248__6_ ( .D(n8366), .CK(clk), .Q(reg_mem[62]) );
  DFF_X1 reg_mem_reg_248__5_ ( .D(n8365), .CK(clk), .Q(reg_mem[61]) );
  DFF_X1 reg_mem_reg_248__4_ ( .D(n8364), .CK(clk), .Q(reg_mem[60]) );
  DFF_X1 reg_mem_reg_248__3_ ( .D(n8363), .CK(clk), .Q(reg_mem[59]) );
  DFF_X1 reg_mem_reg_248__2_ ( .D(n8362), .CK(clk), .Q(reg_mem[58]) );
  DFF_X1 reg_mem_reg_248__1_ ( .D(n8361), .CK(clk), .Q(reg_mem[57]) );
  DFF_X1 reg_mem_reg_248__0_ ( .D(n8360), .CK(clk), .Q(reg_mem[56]) );
  DFF_X1 reg_mem_reg_249__7_ ( .D(n7790), .CK(clk), .Q(reg_mem[55]) );
  DFF_X1 reg_mem_reg_249__6_ ( .D(n7789), .CK(clk), .Q(reg_mem[54]) );
  DFF_X1 reg_mem_reg_249__5_ ( .D(n7788), .CK(clk), .Q(reg_mem[53]) );
  DFF_X1 reg_mem_reg_249__4_ ( .D(n7787), .CK(clk), .Q(reg_mem[52]) );
  DFF_X1 reg_mem_reg_249__3_ ( .D(n7786), .CK(clk), .Q(reg_mem[51]) );
  DFF_X1 reg_mem_reg_249__2_ ( .D(n7785), .CK(clk), .Q(reg_mem[50]) );
  DFF_X1 reg_mem_reg_249__1_ ( .D(n7784), .CK(clk), .Q(reg_mem[49]) );
  DFF_X1 reg_mem_reg_249__0_ ( .D(n7783), .CK(clk), .Q(reg_mem[48]) );
  DFF_X1 reg_mem_reg_250__7_ ( .D(n8943), .CK(clk), .Q(reg_mem[47]) );
  DFF_X1 reg_mem_reg_250__6_ ( .D(n8942), .CK(clk), .Q(reg_mem[46]) );
  DFF_X1 reg_mem_reg_250__5_ ( .D(n8941), .CK(clk), .Q(reg_mem[45]) );
  DFF_X1 reg_mem_reg_250__4_ ( .D(n8940), .CK(clk), .Q(reg_mem[44]) );
  DFF_X1 reg_mem_reg_250__3_ ( .D(n8939), .CK(clk), .Q(reg_mem[43]) );
  DFF_X1 reg_mem_reg_250__2_ ( .D(n8938), .CK(clk), .Q(reg_mem[42]) );
  DFF_X1 reg_mem_reg_250__1_ ( .D(n8937), .CK(clk), .Q(reg_mem[41]) );
  DFF_X1 reg_mem_reg_250__0_ ( .D(n8936), .CK(clk), .Q(reg_mem[40]) );
  DFF_X1 reg_mem_reg_251__7_ ( .D(n7214), .CK(clk), .Q(reg_mem[39]) );
  DFF_X1 reg_mem_reg_251__6_ ( .D(n7213), .CK(clk), .Q(reg_mem[38]) );
  DFF_X1 reg_mem_reg_251__5_ ( .D(n7212), .CK(clk), .Q(reg_mem[37]) );
  DFF_X1 reg_mem_reg_251__4_ ( .D(n7211), .CK(clk), .Q(reg_mem[36]) );
  DFF_X1 reg_mem_reg_251__3_ ( .D(n7210), .CK(clk), .Q(reg_mem[35]) );
  DFF_X1 reg_mem_reg_251__2_ ( .D(n7209), .CK(clk), .Q(reg_mem[34]) );
  DFF_X1 reg_mem_reg_251__1_ ( .D(n7208), .CK(clk), .Q(reg_mem[33]) );
  DFF_X1 reg_mem_reg_251__0_ ( .D(n7207), .CK(clk), .Q(reg_mem[32]) );
  DFF_X1 reg_mem_reg_252__7_ ( .D(n8511), .CK(clk), .Q(reg_mem[31]) );
  DFF_X1 reg_mem_reg_252__6_ ( .D(n8510), .CK(clk), .Q(reg_mem[30]) );
  DFF_X1 reg_mem_reg_252__5_ ( .D(n8509), .CK(clk), .Q(reg_mem[29]) );
  DFF_X1 reg_mem_reg_252__4_ ( .D(n8508), .CK(clk), .Q(reg_mem[28]) );
  DFF_X1 reg_mem_reg_252__3_ ( .D(n8507), .CK(clk), .Q(reg_mem[27]) );
  DFF_X1 reg_mem_reg_252__2_ ( .D(n8506), .CK(clk), .Q(reg_mem[26]) );
  DFF_X1 reg_mem_reg_252__1_ ( .D(n8505), .CK(clk), .Q(reg_mem[25]) );
  DFF_X1 reg_mem_reg_252__0_ ( .D(n8504), .CK(clk), .Q(reg_mem[24]) );
  DFF_X1 reg_mem_reg_253__7_ ( .D(n7934), .CK(clk), .Q(reg_mem[23]) );
  DFF_X1 reg_mem_reg_253__6_ ( .D(n7933), .CK(clk), .Q(reg_mem[22]) );
  DFF_X1 reg_mem_reg_253__5_ ( .D(n7932), .CK(clk), .Q(reg_mem[21]) );
  DFF_X1 reg_mem_reg_253__4_ ( .D(n7931), .CK(clk), .Q(reg_mem[20]) );
  DFF_X1 reg_mem_reg_253__3_ ( .D(n7930), .CK(clk), .Q(reg_mem[19]) );
  DFF_X1 reg_mem_reg_253__2_ ( .D(n7929), .CK(clk), .Q(reg_mem[18]) );
  DFF_X1 reg_mem_reg_253__1_ ( .D(n7928), .CK(clk), .Q(reg_mem[17]) );
  DFF_X1 reg_mem_reg_253__0_ ( .D(n7927), .CK(clk), .Q(reg_mem[16]) );
  DFF_X1 reg_mem_reg_254__7_ ( .D(n9087), .CK(clk), .Q(reg_mem[15]) );
  DFF_X1 reg_mem_reg_254__6_ ( .D(n9086), .CK(clk), .Q(reg_mem[14]) );
  DFF_X1 reg_mem_reg_254__5_ ( .D(n9085), .CK(clk), .Q(reg_mem[13]) );
  DFF_X1 reg_mem_reg_254__4_ ( .D(n9084), .CK(clk), .Q(reg_mem[12]) );
  DFF_X1 reg_mem_reg_254__3_ ( .D(n9083), .CK(clk), .Q(reg_mem[11]) );
  DFF_X1 reg_mem_reg_254__2_ ( .D(n9082), .CK(clk), .Q(reg_mem[10]) );
  DFF_X1 reg_mem_reg_254__1_ ( .D(n9081), .CK(clk), .Q(reg_mem[9]) );
  DFF_X1 reg_mem_reg_254__0_ ( .D(n9080), .CK(clk), .Q(reg_mem[8]) );
  DFF_X1 reg_mem_reg_255__7_ ( .D(n7358), .CK(clk), .Q(reg_mem[7]) );
  DFF_X1 reg_mem_reg_255__6_ ( .D(n7357), .CK(clk), .Q(reg_mem[6]) );
  DFF_X1 reg_mem_reg_255__5_ ( .D(n7356), .CK(clk), .Q(reg_mem[5]) );
  DFF_X1 reg_mem_reg_255__4_ ( .D(n7355), .CK(clk), .Q(reg_mem[4]) );
  DFF_X1 reg_mem_reg_255__3_ ( .D(n7354), .CK(clk), .Q(reg_mem[3]) );
  DFF_X1 reg_mem_reg_255__2_ ( .D(n7353), .CK(clk), .Q(reg_mem[2]) );
  DFF_X1 reg_mem_reg_255__1_ ( .D(n7352), .CK(clk), .Q(reg_mem[1]) );
  DFF_X1 reg_mem_reg_255__0_ ( .D(n7351), .CK(clk), .Q(reg_mem[0]) );
  AND3_X1 U2 ( .A1(n2474), .A2(n2475), .A3(we_s), .ZN(n2323) );
  AND2_X1 U3 ( .A1(n4522), .A2(n4523), .ZN(n2322) );
  AND2_X1 U4 ( .A1(n4533), .A2(n4522), .ZN(n2333) );
  AND2_X1 U5 ( .A1(n4543), .A2(n4522), .ZN(n2343) );
  AND2_X1 U6 ( .A1(n4553), .A2(n4522), .ZN(n2353) );
  AND2_X1 U7 ( .A1(n4563), .A2(n4523), .ZN(n2363) );
  AND2_X1 U8 ( .A1(n4563), .A2(n4533), .ZN(n2373) );
  AND2_X1 U9 ( .A1(n4563), .A2(n4543), .ZN(n2383) );
  AND2_X1 U10 ( .A1(n4563), .A2(n4553), .ZN(n2393) );
  AND2_X1 U11 ( .A1(n4600), .A2(n4523), .ZN(n2403) );
  AND2_X1 U12 ( .A1(n4600), .A2(n4533), .ZN(n2413) );
  AND2_X1 U13 ( .A1(n4600), .A2(n4543), .ZN(n2423) );
  AND2_X1 U14 ( .A1(n4600), .A2(n4553), .ZN(n2433) );
  AND2_X1 U15 ( .A1(n4637), .A2(n4523), .ZN(n2443) );
  AND2_X1 U16 ( .A1(n4637), .A2(n4533), .ZN(n2453) );
  AND2_X1 U17 ( .A1(n4637), .A2(n4543), .ZN(n2463) );
  AND2_X1 U18 ( .A1(n4637), .A2(n4553), .ZN(n2473) );
  INV_X1 U19 ( .A(n2314), .ZN(n7359) );
  INV_X1 U20 ( .A(n2915), .ZN(n7323) );
  INV_X1 U21 ( .A(n2925), .ZN(n9052) );
  INV_X1 U22 ( .A(n2934), .ZN(n7899) );
  INV_X1 U23 ( .A(n2943), .ZN(n8476) );
  INV_X1 U24 ( .A(n2952), .ZN(n7179) );
  INV_X1 U25 ( .A(n2961), .ZN(n8908) );
  INV_X1 U26 ( .A(n2970), .ZN(n7755) );
  INV_X1 U27 ( .A(n2979), .ZN(n8332) );
  INV_X1 U28 ( .A(n2988), .ZN(n7035) );
  INV_X1 U29 ( .A(n2997), .ZN(n8764) );
  INV_X1 U30 ( .A(n3006), .ZN(n7611) );
  INV_X1 U31 ( .A(n3015), .ZN(n8188) );
  INV_X1 U32 ( .A(n3024), .ZN(n6891) );
  INV_X1 U33 ( .A(n3033), .ZN(n8620) );
  INV_X1 U34 ( .A(n3042), .ZN(n7467) );
  INV_X1 U35 ( .A(n3051), .ZN(n8044) );
  INV_X1 U36 ( .A(n3061), .ZN(n7314) );
  INV_X1 U37 ( .A(n3071), .ZN(n9043) );
  INV_X1 U38 ( .A(n3080), .ZN(n7890) );
  INV_X1 U39 ( .A(n3089), .ZN(n8467) );
  INV_X1 U40 ( .A(n3098), .ZN(n7170) );
  INV_X1 U41 ( .A(n3107), .ZN(n8899) );
  INV_X1 U42 ( .A(n3116), .ZN(n7746) );
  INV_X1 U43 ( .A(n3125), .ZN(n8323) );
  INV_X1 U44 ( .A(n3134), .ZN(n7026) );
  INV_X1 U45 ( .A(n3143), .ZN(n8755) );
  INV_X1 U46 ( .A(n3152), .ZN(n7602) );
  INV_X1 U47 ( .A(n3161), .ZN(n8179) );
  INV_X1 U48 ( .A(n3170), .ZN(n6882) );
  INV_X1 U49 ( .A(n3179), .ZN(n8611) );
  INV_X1 U50 ( .A(n3188), .ZN(n7458) );
  INV_X1 U51 ( .A(n3197), .ZN(n8035) );
  INV_X1 U52 ( .A(n3206), .ZN(n7305) );
  INV_X1 U53 ( .A(n3216), .ZN(n9034) );
  INV_X1 U54 ( .A(n3225), .ZN(n7881) );
  INV_X1 U55 ( .A(n3234), .ZN(n8458) );
  INV_X1 U56 ( .A(n3243), .ZN(n7161) );
  INV_X1 U57 ( .A(n3252), .ZN(n8890) );
  INV_X1 U58 ( .A(n3261), .ZN(n7737) );
  INV_X1 U59 ( .A(n3270), .ZN(n8314) );
  INV_X1 U60 ( .A(n3279), .ZN(n7017) );
  INV_X1 U61 ( .A(n3288), .ZN(n8746) );
  INV_X1 U62 ( .A(n3297), .ZN(n7593) );
  INV_X1 U63 ( .A(n3306), .ZN(n8170) );
  INV_X1 U64 ( .A(n3315), .ZN(n6873) );
  INV_X1 U65 ( .A(n3324), .ZN(n8602) );
  INV_X1 U66 ( .A(n3333), .ZN(n7449) );
  INV_X1 U67 ( .A(n3342), .ZN(n8026) );
  INV_X1 U68 ( .A(n3351), .ZN(n7296) );
  INV_X1 U69 ( .A(n3361), .ZN(n9025) );
  INV_X1 U70 ( .A(n3370), .ZN(n7872) );
  INV_X1 U71 ( .A(n3379), .ZN(n8449) );
  INV_X1 U72 ( .A(n3388), .ZN(n7152) );
  INV_X1 U73 ( .A(n3397), .ZN(n8881) );
  INV_X1 U74 ( .A(n3406), .ZN(n7728) );
  INV_X1 U75 ( .A(n3415), .ZN(n8305) );
  INV_X1 U76 ( .A(n3424), .ZN(n7008) );
  INV_X1 U77 ( .A(n3433), .ZN(n8737) );
  INV_X1 U78 ( .A(n3442), .ZN(n7584) );
  INV_X1 U79 ( .A(n3451), .ZN(n8161) );
  INV_X1 U80 ( .A(n3460), .ZN(n6864) );
  INV_X1 U81 ( .A(n3469), .ZN(n8593) );
  INV_X1 U82 ( .A(n3478), .ZN(n7440) );
  INV_X1 U83 ( .A(n3487), .ZN(n8017) );
  INV_X1 U84 ( .A(n3496), .ZN(n7287) );
  INV_X1 U85 ( .A(n3506), .ZN(n9016) );
  INV_X1 U86 ( .A(n3515), .ZN(n7863) );
  INV_X1 U87 ( .A(n3524), .ZN(n8440) );
  INV_X1 U88 ( .A(n3533), .ZN(n7143) );
  INV_X1 U89 ( .A(n3542), .ZN(n8872) );
  INV_X1 U90 ( .A(n3551), .ZN(n7719) );
  INV_X1 U91 ( .A(n3560), .ZN(n8296) );
  INV_X1 U92 ( .A(n3569), .ZN(n6999) );
  INV_X1 U93 ( .A(n3578), .ZN(n8728) );
  INV_X1 U94 ( .A(n3587), .ZN(n7575) );
  INV_X1 U95 ( .A(n3596), .ZN(n8152) );
  INV_X1 U96 ( .A(n3605), .ZN(n6855) );
  INV_X1 U97 ( .A(n3614), .ZN(n8584) );
  INV_X1 U98 ( .A(n3623), .ZN(n7431) );
  INV_X1 U99 ( .A(n3632), .ZN(n8008) );
  INV_X1 U100 ( .A(n3642), .ZN(n7278) );
  INV_X1 U101 ( .A(n3652), .ZN(n9007) );
  INV_X1 U102 ( .A(n3661), .ZN(n7854) );
  INV_X1 U103 ( .A(n3670), .ZN(n8431) );
  INV_X1 U104 ( .A(n3679), .ZN(n7134) );
  INV_X1 U105 ( .A(n3688), .ZN(n8863) );
  INV_X1 U106 ( .A(n3697), .ZN(n7710) );
  INV_X1 U107 ( .A(n3706), .ZN(n8287) );
  INV_X1 U108 ( .A(n3715), .ZN(n6990) );
  INV_X1 U109 ( .A(n3724), .ZN(n8719) );
  INV_X1 U110 ( .A(n3733), .ZN(n7566) );
  INV_X1 U111 ( .A(n3742), .ZN(n8143) );
  INV_X1 U112 ( .A(n3751), .ZN(n6846) );
  INV_X1 U113 ( .A(n3760), .ZN(n8575) );
  INV_X1 U114 ( .A(n3769), .ZN(n7422) );
  INV_X1 U115 ( .A(n3778), .ZN(n7999) );
  INV_X1 U116 ( .A(n3787), .ZN(n7269) );
  INV_X1 U117 ( .A(n3797), .ZN(n8998) );
  INV_X1 U118 ( .A(n3806), .ZN(n7845) );
  INV_X1 U119 ( .A(n3815), .ZN(n8422) );
  INV_X1 U120 ( .A(n3824), .ZN(n7125) );
  INV_X1 U121 ( .A(n3833), .ZN(n8854) );
  INV_X1 U122 ( .A(n3842), .ZN(n7701) );
  INV_X1 U123 ( .A(n3851), .ZN(n8278) );
  INV_X1 U124 ( .A(n3860), .ZN(n6981) );
  INV_X1 U125 ( .A(n3869), .ZN(n8710) );
  INV_X1 U126 ( .A(n3878), .ZN(n7557) );
  INV_X1 U127 ( .A(n3887), .ZN(n8134) );
  INV_X1 U128 ( .A(n3896), .ZN(n6837) );
  INV_X1 U129 ( .A(n3905), .ZN(n8566) );
  INV_X1 U130 ( .A(n3914), .ZN(n7413) );
  INV_X1 U131 ( .A(n3923), .ZN(n7990) );
  INV_X1 U132 ( .A(n3932), .ZN(n7260) );
  INV_X1 U133 ( .A(n3942), .ZN(n8989) );
  INV_X1 U134 ( .A(n3951), .ZN(n7836) );
  INV_X1 U135 ( .A(n3960), .ZN(n8413) );
  INV_X1 U136 ( .A(n3969), .ZN(n7116) );
  INV_X1 U137 ( .A(n3978), .ZN(n8845) );
  INV_X1 U138 ( .A(n3987), .ZN(n7692) );
  INV_X1 U139 ( .A(n3996), .ZN(n8269) );
  INV_X1 U140 ( .A(n4005), .ZN(n6972) );
  INV_X1 U141 ( .A(n4014), .ZN(n8701) );
  INV_X1 U142 ( .A(n4023), .ZN(n7548) );
  INV_X1 U143 ( .A(n4032), .ZN(n8125) );
  INV_X1 U144 ( .A(n4041), .ZN(n6828) );
  INV_X1 U145 ( .A(n4050), .ZN(n8557) );
  INV_X1 U146 ( .A(n4059), .ZN(n7404) );
  INV_X1 U147 ( .A(n4068), .ZN(n7981) );
  INV_X1 U148 ( .A(n4223), .ZN(n7242) );
  INV_X1 U149 ( .A(n4233), .ZN(n8971) );
  INV_X1 U150 ( .A(n4242), .ZN(n7818) );
  INV_X1 U151 ( .A(n4251), .ZN(n8395) );
  INV_X1 U152 ( .A(n4260), .ZN(n7098) );
  INV_X1 U153 ( .A(n4269), .ZN(n8827) );
  INV_X1 U154 ( .A(n4278), .ZN(n7674) );
  INV_X1 U155 ( .A(n4287), .ZN(n8251) );
  INV_X1 U156 ( .A(n4296), .ZN(n6954) );
  INV_X1 U157 ( .A(n4305), .ZN(n8683) );
  INV_X1 U158 ( .A(n4314), .ZN(n7530) );
  INV_X1 U159 ( .A(n4323), .ZN(n8107) );
  INV_X1 U160 ( .A(n4332), .ZN(n6810) );
  INV_X1 U161 ( .A(n4341), .ZN(n8539) );
  INV_X1 U162 ( .A(n4350), .ZN(n7386) );
  INV_X1 U163 ( .A(n4359), .ZN(n7963) );
  INV_X1 U164 ( .A(n4368), .ZN(n7233) );
  INV_X1 U165 ( .A(n4378), .ZN(n8962) );
  INV_X1 U166 ( .A(n4387), .ZN(n7809) );
  INV_X1 U167 ( .A(n4396), .ZN(n8386) );
  INV_X1 U168 ( .A(n4405), .ZN(n7089) );
  INV_X1 U169 ( .A(n4414), .ZN(n8818) );
  INV_X1 U170 ( .A(n4423), .ZN(n7665) );
  INV_X1 U171 ( .A(n4432), .ZN(n8242) );
  INV_X1 U172 ( .A(n4441), .ZN(n6945) );
  INV_X1 U173 ( .A(n4450), .ZN(n8674) );
  INV_X1 U174 ( .A(n4459), .ZN(n7521) );
  INV_X1 U175 ( .A(n4468), .ZN(n8098) );
  INV_X1 U176 ( .A(n4477), .ZN(n6801) );
  INV_X1 U177 ( .A(n4486), .ZN(n8530) );
  INV_X1 U178 ( .A(n4495), .ZN(n7377) );
  INV_X1 U179 ( .A(n4504), .ZN(n7954) );
  INV_X1 U180 ( .A(n4513), .ZN(n7224) );
  INV_X1 U181 ( .A(n4525), .ZN(n8953) );
  INV_X1 U182 ( .A(n4535), .ZN(n7800) );
  INV_X1 U183 ( .A(n4545), .ZN(n8377) );
  INV_X1 U184 ( .A(n4555), .ZN(n7080) );
  INV_X1 U185 ( .A(n4565), .ZN(n8809) );
  INV_X1 U186 ( .A(n4574), .ZN(n7656) );
  INV_X1 U187 ( .A(n4583), .ZN(n8233) );
  INV_X1 U188 ( .A(n4592), .ZN(n6936) );
  INV_X1 U189 ( .A(n4602), .ZN(n8665) );
  INV_X1 U190 ( .A(n4611), .ZN(n7512) );
  INV_X1 U191 ( .A(n4620), .ZN(n8089) );
  INV_X1 U192 ( .A(n4629), .ZN(n6792) );
  INV_X1 U193 ( .A(n4639), .ZN(n8521) );
  INV_X1 U194 ( .A(n4648), .ZN(n7368) );
  INV_X1 U195 ( .A(n4657), .ZN(n7945) );
  INV_X1 U196 ( .A(n2325), .ZN(n9088) );
  INV_X1 U197 ( .A(n2335), .ZN(n7935) );
  INV_X1 U198 ( .A(n2345), .ZN(n8512) );
  INV_X1 U199 ( .A(n2355), .ZN(n7215) );
  INV_X1 U200 ( .A(n2365), .ZN(n8944) );
  INV_X1 U201 ( .A(n2375), .ZN(n7791) );
  INV_X1 U202 ( .A(n2385), .ZN(n8368) );
  INV_X1 U203 ( .A(n2395), .ZN(n7071) );
  INV_X1 U204 ( .A(n2405), .ZN(n8800) );
  INV_X1 U205 ( .A(n2415), .ZN(n7647) );
  INV_X1 U206 ( .A(n2425), .ZN(n8224) );
  INV_X1 U207 ( .A(n2435), .ZN(n6927) );
  INV_X1 U208 ( .A(n2445), .ZN(n8656) );
  INV_X1 U209 ( .A(n2455), .ZN(n7503) );
  INV_X1 U210 ( .A(n2465), .ZN(n8080) );
  INV_X1 U211 ( .A(n2477), .ZN(n7350) );
  INV_X1 U212 ( .A(n2487), .ZN(n9079) );
  INV_X1 U213 ( .A(n2496), .ZN(n7926) );
  INV_X1 U214 ( .A(n2505), .ZN(n8503) );
  INV_X1 U215 ( .A(n2514), .ZN(n7206) );
  INV_X1 U216 ( .A(n2523), .ZN(n8935) );
  INV_X1 U217 ( .A(n2532), .ZN(n7782) );
  INV_X1 U218 ( .A(n2541), .ZN(n8359) );
  INV_X1 U219 ( .A(n2550), .ZN(n7062) );
  INV_X1 U220 ( .A(n2559), .ZN(n8791) );
  INV_X1 U221 ( .A(n2568), .ZN(n7638) );
  INV_X1 U222 ( .A(n2577), .ZN(n8215) );
  INV_X1 U223 ( .A(n2586), .ZN(n6918) );
  INV_X1 U224 ( .A(n2595), .ZN(n8647) );
  INV_X1 U225 ( .A(n2604), .ZN(n7494) );
  INV_X1 U226 ( .A(n2613), .ZN(n8071) );
  INV_X1 U227 ( .A(n2623), .ZN(n7341) );
  INV_X1 U228 ( .A(n2633), .ZN(n9070) );
  INV_X1 U229 ( .A(n2642), .ZN(n7917) );
  INV_X1 U230 ( .A(n2651), .ZN(n8494) );
  INV_X1 U231 ( .A(n2660), .ZN(n7197) );
  INV_X1 U232 ( .A(n2669), .ZN(n8926) );
  INV_X1 U233 ( .A(n2678), .ZN(n7773) );
  INV_X1 U234 ( .A(n2687), .ZN(n8350) );
  INV_X1 U235 ( .A(n2696), .ZN(n7053) );
  INV_X1 U236 ( .A(n2705), .ZN(n8782) );
  INV_X1 U237 ( .A(n2714), .ZN(n7629) );
  INV_X1 U238 ( .A(n2723), .ZN(n8206) );
  INV_X1 U239 ( .A(n2732), .ZN(n6909) );
  INV_X1 U240 ( .A(n2741), .ZN(n8638) );
  INV_X1 U241 ( .A(n2750), .ZN(n7485) );
  INV_X1 U242 ( .A(n2759), .ZN(n8062) );
  INV_X1 U243 ( .A(n2769), .ZN(n7332) );
  INV_X1 U244 ( .A(n2779), .ZN(n9061) );
  INV_X1 U245 ( .A(n2788), .ZN(n7908) );
  INV_X1 U246 ( .A(n2797), .ZN(n8485) );
  INV_X1 U247 ( .A(n2806), .ZN(n7188) );
  INV_X1 U248 ( .A(n2815), .ZN(n8917) );
  INV_X1 U249 ( .A(n2824), .ZN(n7764) );
  INV_X1 U250 ( .A(n2833), .ZN(n8341) );
  INV_X1 U251 ( .A(n2842), .ZN(n7044) );
  INV_X1 U252 ( .A(n2851), .ZN(n8773) );
  INV_X1 U253 ( .A(n2860), .ZN(n7620) );
  INV_X1 U254 ( .A(n2869), .ZN(n8197) );
  INV_X1 U255 ( .A(n2878), .ZN(n6900) );
  INV_X1 U256 ( .A(n2887), .ZN(n8629) );
  INV_X1 U257 ( .A(n2896), .ZN(n7476) );
  INV_X1 U258 ( .A(n2905), .ZN(n8053) );
  INV_X1 U259 ( .A(n4077), .ZN(n7251) );
  INV_X1 U260 ( .A(n4087), .ZN(n8980) );
  INV_X1 U261 ( .A(n4096), .ZN(n7827) );
  INV_X1 U262 ( .A(n4105), .ZN(n8404) );
  INV_X1 U263 ( .A(n4114), .ZN(n7107) );
  INV_X1 U264 ( .A(n4123), .ZN(n8836) );
  INV_X1 U265 ( .A(n4132), .ZN(n7683) );
  INV_X1 U266 ( .A(n4141), .ZN(n8260) );
  INV_X1 U267 ( .A(n4150), .ZN(n6963) );
  INV_X1 U268 ( .A(n4159), .ZN(n8692) );
  INV_X1 U269 ( .A(n4168), .ZN(n7539) );
  INV_X1 U270 ( .A(n4177), .ZN(n8116) );
  INV_X1 U271 ( .A(n4186), .ZN(n6819) );
  INV_X1 U272 ( .A(n4195), .ZN(n8548) );
  INV_X1 U273 ( .A(n4204), .ZN(n7395) );
  INV_X1 U274 ( .A(n4213), .ZN(n7972) );
  NAND2_X1 U275 ( .A1(n2923), .A2(n2322), .ZN(n2915) );
  NAND2_X1 U276 ( .A1(n2923), .A2(n2333), .ZN(n2925) );
  NAND2_X1 U277 ( .A1(n2923), .A2(n2343), .ZN(n2934) );
  NAND2_X1 U278 ( .A1(n2923), .A2(n2353), .ZN(n2943) );
  NAND2_X1 U279 ( .A1(n2923), .A2(n2363), .ZN(n2952) );
  NAND2_X1 U280 ( .A1(n2923), .A2(n2373), .ZN(n2961) );
  NAND2_X1 U281 ( .A1(n2923), .A2(n2383), .ZN(n2970) );
  NAND2_X1 U282 ( .A1(n2923), .A2(n2393), .ZN(n2979) );
  NAND2_X1 U283 ( .A1(n2923), .A2(n2403), .ZN(n2988) );
  NAND2_X1 U284 ( .A1(n2923), .A2(n2413), .ZN(n2997) );
  NAND2_X1 U285 ( .A1(n2923), .A2(n2423), .ZN(n3006) );
  NAND2_X1 U286 ( .A1(n2923), .A2(n2433), .ZN(n3015) );
  NAND2_X1 U287 ( .A1(n2923), .A2(n2443), .ZN(n3024) );
  NAND2_X1 U288 ( .A1(n2923), .A2(n2453), .ZN(n3033) );
  NAND2_X1 U289 ( .A1(n2923), .A2(n2463), .ZN(n3042) );
  NAND2_X1 U290 ( .A1(n2923), .A2(n2473), .ZN(n3051) );
  NAND2_X1 U291 ( .A1(n3069), .A2(n2322), .ZN(n3061) );
  NAND2_X1 U292 ( .A1(n3069), .A2(n2333), .ZN(n3071) );
  NAND2_X1 U293 ( .A1(n3069), .A2(n2343), .ZN(n3080) );
  NAND2_X1 U294 ( .A1(n3069), .A2(n2353), .ZN(n3089) );
  NAND2_X1 U295 ( .A1(n3069), .A2(n2363), .ZN(n3098) );
  NAND2_X1 U296 ( .A1(n3069), .A2(n2373), .ZN(n3107) );
  NAND2_X1 U297 ( .A1(n3069), .A2(n2383), .ZN(n3116) );
  NAND2_X1 U298 ( .A1(n3069), .A2(n2393), .ZN(n3125) );
  NAND2_X1 U299 ( .A1(n3069), .A2(n2403), .ZN(n3134) );
  NAND2_X1 U300 ( .A1(n3069), .A2(n2413), .ZN(n3143) );
  NAND2_X1 U301 ( .A1(n3069), .A2(n2423), .ZN(n3152) );
  NAND2_X1 U302 ( .A1(n3069), .A2(n2433), .ZN(n3161) );
  NAND2_X1 U303 ( .A1(n3069), .A2(n2443), .ZN(n3170) );
  NAND2_X1 U304 ( .A1(n3069), .A2(n2453), .ZN(n3179) );
  NAND2_X1 U305 ( .A1(n3069), .A2(n2463), .ZN(n3188) );
  NAND2_X1 U306 ( .A1(n3069), .A2(n2473), .ZN(n3197) );
  NAND2_X1 U307 ( .A1(n3214), .A2(n2322), .ZN(n3206) );
  NAND2_X1 U308 ( .A1(n3214), .A2(n2333), .ZN(n3216) );
  NAND2_X1 U309 ( .A1(n3214), .A2(n2343), .ZN(n3225) );
  NAND2_X1 U310 ( .A1(n3214), .A2(n2353), .ZN(n3234) );
  NAND2_X1 U311 ( .A1(n3214), .A2(n2363), .ZN(n3243) );
  NAND2_X1 U312 ( .A1(n3214), .A2(n2373), .ZN(n3252) );
  NAND2_X1 U313 ( .A1(n3214), .A2(n2383), .ZN(n3261) );
  NAND2_X1 U314 ( .A1(n3214), .A2(n2393), .ZN(n3270) );
  NAND2_X1 U315 ( .A1(n3214), .A2(n2403), .ZN(n3279) );
  NAND2_X1 U316 ( .A1(n3214), .A2(n2413), .ZN(n3288) );
  NAND2_X1 U317 ( .A1(n3214), .A2(n2423), .ZN(n3297) );
  NAND2_X1 U318 ( .A1(n3214), .A2(n2433), .ZN(n3306) );
  NAND2_X1 U319 ( .A1(n3214), .A2(n2443), .ZN(n3315) );
  NAND2_X1 U320 ( .A1(n3214), .A2(n2453), .ZN(n3324) );
  NAND2_X1 U321 ( .A1(n3214), .A2(n2463), .ZN(n3333) );
  NAND2_X1 U322 ( .A1(n3214), .A2(n2473), .ZN(n3342) );
  NAND2_X1 U323 ( .A1(n3359), .A2(n2322), .ZN(n3351) );
  NAND2_X1 U324 ( .A1(n3359), .A2(n2333), .ZN(n3361) );
  NAND2_X1 U325 ( .A1(n3359), .A2(n2343), .ZN(n3370) );
  NAND2_X1 U326 ( .A1(n3359), .A2(n2353), .ZN(n3379) );
  NAND2_X1 U327 ( .A1(n3359), .A2(n2363), .ZN(n3388) );
  NAND2_X1 U328 ( .A1(n3359), .A2(n2373), .ZN(n3397) );
  NAND2_X1 U329 ( .A1(n3359), .A2(n2383), .ZN(n3406) );
  NAND2_X1 U330 ( .A1(n3359), .A2(n2393), .ZN(n3415) );
  NAND2_X1 U331 ( .A1(n3359), .A2(n2403), .ZN(n3424) );
  NAND2_X1 U332 ( .A1(n3359), .A2(n2413), .ZN(n3433) );
  NAND2_X1 U333 ( .A1(n3359), .A2(n2423), .ZN(n3442) );
  NAND2_X1 U334 ( .A1(n3359), .A2(n2433), .ZN(n3451) );
  NAND2_X1 U335 ( .A1(n3359), .A2(n2443), .ZN(n3460) );
  NAND2_X1 U336 ( .A1(n3359), .A2(n2453), .ZN(n3469) );
  NAND2_X1 U337 ( .A1(n3359), .A2(n2463), .ZN(n3478) );
  NAND2_X1 U338 ( .A1(n3359), .A2(n2473), .ZN(n3487) );
  NAND2_X1 U339 ( .A1(n3504), .A2(n2322), .ZN(n3496) );
  NAND2_X1 U340 ( .A1(n3504), .A2(n2333), .ZN(n3506) );
  NAND2_X1 U341 ( .A1(n3504), .A2(n2343), .ZN(n3515) );
  NAND2_X1 U342 ( .A1(n3504), .A2(n2353), .ZN(n3524) );
  NAND2_X1 U343 ( .A1(n3504), .A2(n2363), .ZN(n3533) );
  NAND2_X1 U344 ( .A1(n3504), .A2(n2373), .ZN(n3542) );
  NAND2_X1 U345 ( .A1(n3504), .A2(n2383), .ZN(n3551) );
  NAND2_X1 U346 ( .A1(n3504), .A2(n2393), .ZN(n3560) );
  NAND2_X1 U347 ( .A1(n3504), .A2(n2403), .ZN(n3569) );
  NAND2_X1 U348 ( .A1(n3504), .A2(n2413), .ZN(n3578) );
  NAND2_X1 U349 ( .A1(n3504), .A2(n2423), .ZN(n3587) );
  NAND2_X1 U350 ( .A1(n3504), .A2(n2433), .ZN(n3596) );
  NAND2_X1 U351 ( .A1(n3504), .A2(n2443), .ZN(n3605) );
  NAND2_X1 U352 ( .A1(n3504), .A2(n2453), .ZN(n3614) );
  NAND2_X1 U353 ( .A1(n3504), .A2(n2463), .ZN(n3623) );
  NAND2_X1 U354 ( .A1(n3504), .A2(n2473), .ZN(n3632) );
  NAND2_X1 U355 ( .A1(n3650), .A2(n2322), .ZN(n3642) );
  NAND2_X1 U356 ( .A1(n3650), .A2(n2333), .ZN(n3652) );
  NAND2_X1 U357 ( .A1(n3650), .A2(n2343), .ZN(n3661) );
  NAND2_X1 U358 ( .A1(n3650), .A2(n2353), .ZN(n3670) );
  NAND2_X1 U359 ( .A1(n3650), .A2(n2363), .ZN(n3679) );
  NAND2_X1 U360 ( .A1(n3650), .A2(n2373), .ZN(n3688) );
  NAND2_X1 U361 ( .A1(n3650), .A2(n2383), .ZN(n3697) );
  NAND2_X1 U362 ( .A1(n3650), .A2(n2393), .ZN(n3706) );
  NAND2_X1 U363 ( .A1(n3650), .A2(n2403), .ZN(n3715) );
  NAND2_X1 U364 ( .A1(n3650), .A2(n2413), .ZN(n3724) );
  NAND2_X1 U365 ( .A1(n3650), .A2(n2423), .ZN(n3733) );
  NAND2_X1 U366 ( .A1(n3650), .A2(n2433), .ZN(n3742) );
  NAND2_X1 U367 ( .A1(n3650), .A2(n2443), .ZN(n3751) );
  NAND2_X1 U368 ( .A1(n3650), .A2(n2453), .ZN(n3760) );
  NAND2_X1 U369 ( .A1(n3650), .A2(n2463), .ZN(n3769) );
  NAND2_X1 U370 ( .A1(n3650), .A2(n2473), .ZN(n3778) );
  NAND2_X1 U371 ( .A1(n3795), .A2(n2322), .ZN(n3787) );
  NAND2_X1 U372 ( .A1(n3795), .A2(n2333), .ZN(n3797) );
  NAND2_X1 U373 ( .A1(n3795), .A2(n2343), .ZN(n3806) );
  NAND2_X1 U374 ( .A1(n3795), .A2(n2353), .ZN(n3815) );
  NAND2_X1 U375 ( .A1(n3795), .A2(n2363), .ZN(n3824) );
  NAND2_X1 U376 ( .A1(n3795), .A2(n2373), .ZN(n3833) );
  NAND2_X1 U377 ( .A1(n3795), .A2(n2383), .ZN(n3842) );
  NAND2_X1 U378 ( .A1(n3795), .A2(n2393), .ZN(n3851) );
  NAND2_X1 U379 ( .A1(n3795), .A2(n2403), .ZN(n3860) );
  NAND2_X1 U380 ( .A1(n3795), .A2(n2413), .ZN(n3869) );
  NAND2_X1 U381 ( .A1(n3795), .A2(n2423), .ZN(n3878) );
  NAND2_X1 U382 ( .A1(n3795), .A2(n2433), .ZN(n3887) );
  NAND2_X1 U383 ( .A1(n3795), .A2(n2443), .ZN(n3896) );
  NAND2_X1 U384 ( .A1(n3795), .A2(n2453), .ZN(n3905) );
  NAND2_X1 U385 ( .A1(n3795), .A2(n2463), .ZN(n3914) );
  NAND2_X1 U386 ( .A1(n3795), .A2(n2473), .ZN(n3923) );
  NAND2_X1 U387 ( .A1(n3940), .A2(n2322), .ZN(n3932) );
  NAND2_X1 U388 ( .A1(n3940), .A2(n2333), .ZN(n3942) );
  NAND2_X1 U389 ( .A1(n3940), .A2(n2343), .ZN(n3951) );
  NAND2_X1 U390 ( .A1(n3940), .A2(n2353), .ZN(n3960) );
  NAND2_X1 U391 ( .A1(n3940), .A2(n2363), .ZN(n3969) );
  NAND2_X1 U392 ( .A1(n3940), .A2(n2373), .ZN(n3978) );
  NAND2_X1 U393 ( .A1(n3940), .A2(n2383), .ZN(n3987) );
  NAND2_X1 U394 ( .A1(n3940), .A2(n2393), .ZN(n3996) );
  NAND2_X1 U395 ( .A1(n3940), .A2(n2403), .ZN(n4005) );
  NAND2_X1 U396 ( .A1(n3940), .A2(n2413), .ZN(n4014) );
  NAND2_X1 U397 ( .A1(n3940), .A2(n2423), .ZN(n4023) );
  NAND2_X1 U398 ( .A1(n3940), .A2(n2433), .ZN(n4032) );
  NAND2_X1 U399 ( .A1(n3940), .A2(n2443), .ZN(n4041) );
  NAND2_X1 U400 ( .A1(n3940), .A2(n2453), .ZN(n4050) );
  NAND2_X1 U401 ( .A1(n3940), .A2(n2463), .ZN(n4059) );
  NAND2_X1 U402 ( .A1(n3940), .A2(n2473), .ZN(n4068) );
  NAND2_X1 U403 ( .A1(n4231), .A2(n2322), .ZN(n4223) );
  NAND2_X1 U404 ( .A1(n4231), .A2(n2333), .ZN(n4233) );
  NAND2_X1 U405 ( .A1(n4231), .A2(n2343), .ZN(n4242) );
  NAND2_X1 U406 ( .A1(n4231), .A2(n2353), .ZN(n4251) );
  NAND2_X1 U407 ( .A1(n4231), .A2(n2363), .ZN(n4260) );
  NAND2_X1 U408 ( .A1(n4231), .A2(n2373), .ZN(n4269) );
  NAND2_X1 U409 ( .A1(n4231), .A2(n2383), .ZN(n4278) );
  NAND2_X1 U410 ( .A1(n4231), .A2(n2393), .ZN(n4287) );
  NAND2_X1 U411 ( .A1(n4231), .A2(n2403), .ZN(n4296) );
  NAND2_X1 U412 ( .A1(n4231), .A2(n2413), .ZN(n4305) );
  NAND2_X1 U413 ( .A1(n4231), .A2(n2423), .ZN(n4314) );
  NAND2_X1 U414 ( .A1(n4231), .A2(n2433), .ZN(n4323) );
  NAND2_X1 U415 ( .A1(n4231), .A2(n2443), .ZN(n4332) );
  NAND2_X1 U416 ( .A1(n4231), .A2(n2453), .ZN(n4341) );
  NAND2_X1 U417 ( .A1(n4231), .A2(n2463), .ZN(n4350) );
  NAND2_X1 U418 ( .A1(n4231), .A2(n2473), .ZN(n4359) );
  NAND2_X1 U419 ( .A1(n4376), .A2(n2322), .ZN(n4368) );
  NAND2_X1 U420 ( .A1(n4376), .A2(n2333), .ZN(n4378) );
  NAND2_X1 U421 ( .A1(n4376), .A2(n2343), .ZN(n4387) );
  NAND2_X1 U422 ( .A1(n4376), .A2(n2353), .ZN(n4396) );
  NAND2_X1 U423 ( .A1(n4376), .A2(n2363), .ZN(n4405) );
  NAND2_X1 U424 ( .A1(n4376), .A2(n2373), .ZN(n4414) );
  NAND2_X1 U425 ( .A1(n4376), .A2(n2383), .ZN(n4423) );
  NAND2_X1 U426 ( .A1(n4376), .A2(n2393), .ZN(n4432) );
  NAND2_X1 U427 ( .A1(n4376), .A2(n2403), .ZN(n4441) );
  NAND2_X1 U428 ( .A1(n4376), .A2(n2413), .ZN(n4450) );
  NAND2_X1 U429 ( .A1(n4376), .A2(n2423), .ZN(n4459) );
  NAND2_X1 U430 ( .A1(n4376), .A2(n2433), .ZN(n4468) );
  NAND2_X1 U431 ( .A1(n4376), .A2(n2443), .ZN(n4477) );
  NAND2_X1 U432 ( .A1(n4376), .A2(n2453), .ZN(n4486) );
  NAND2_X1 U433 ( .A1(n4376), .A2(n2463), .ZN(n4495) );
  NAND2_X1 U434 ( .A1(n4376), .A2(n2473), .ZN(n4504) );
  NAND2_X1 U435 ( .A1(n4521), .A2(n2322), .ZN(n4513) );
  NAND2_X1 U436 ( .A1(n4521), .A2(n2333), .ZN(n4525) );
  NAND2_X1 U437 ( .A1(n4521), .A2(n2343), .ZN(n4535) );
  NAND2_X1 U438 ( .A1(n4521), .A2(n2353), .ZN(n4545) );
  NAND2_X1 U439 ( .A1(n4521), .A2(n2363), .ZN(n4555) );
  NAND2_X1 U440 ( .A1(n4521), .A2(n2373), .ZN(n4565) );
  NAND2_X1 U441 ( .A1(n4521), .A2(n2383), .ZN(n4574) );
  NAND2_X1 U442 ( .A1(n4521), .A2(n2393), .ZN(n4583) );
  NAND2_X1 U443 ( .A1(n4521), .A2(n2403), .ZN(n4592) );
  NAND2_X1 U444 ( .A1(n4521), .A2(n2413), .ZN(n4602) );
  NAND2_X1 U445 ( .A1(n4521), .A2(n2423), .ZN(n4611) );
  NAND2_X1 U446 ( .A1(n4521), .A2(n2433), .ZN(n4620) );
  NAND2_X1 U447 ( .A1(n4521), .A2(n2443), .ZN(n4629) );
  NAND2_X1 U448 ( .A1(n4521), .A2(n2453), .ZN(n4639) );
  NAND2_X1 U449 ( .A1(n4521), .A2(n2463), .ZN(n4648) );
  NAND2_X1 U450 ( .A1(n4521), .A2(n2473), .ZN(n4657) );
  NAND2_X1 U451 ( .A1(n2322), .A2(n2323), .ZN(n2314) );
  NAND2_X1 U452 ( .A1(n2333), .A2(n2323), .ZN(n2325) );
  NAND2_X1 U453 ( .A1(n2343), .A2(n2323), .ZN(n2335) );
  NAND2_X1 U454 ( .A1(n2353), .A2(n2323), .ZN(n2345) );
  NAND2_X1 U455 ( .A1(n2363), .A2(n2323), .ZN(n2355) );
  NAND2_X1 U456 ( .A1(n2373), .A2(n2323), .ZN(n2365) );
  NAND2_X1 U457 ( .A1(n2383), .A2(n2323), .ZN(n2375) );
  NAND2_X1 U458 ( .A1(n2393), .A2(n2323), .ZN(n2385) );
  NAND2_X1 U459 ( .A1(n2403), .A2(n2323), .ZN(n2395) );
  NAND2_X1 U460 ( .A1(n2413), .A2(n2323), .ZN(n2405) );
  NAND2_X1 U461 ( .A1(n2423), .A2(n2323), .ZN(n2415) );
  NAND2_X1 U462 ( .A1(n2433), .A2(n2323), .ZN(n2425) );
  NAND2_X1 U463 ( .A1(n2443), .A2(n2323), .ZN(n2435) );
  NAND2_X1 U464 ( .A1(n2453), .A2(n2323), .ZN(n2445) );
  NAND2_X1 U465 ( .A1(n2463), .A2(n2323), .ZN(n2455) );
  NAND2_X1 U466 ( .A1(n2473), .A2(n2323), .ZN(n2465) );
  NAND2_X1 U467 ( .A1(n2485), .A2(n2322), .ZN(n2477) );
  NAND2_X1 U468 ( .A1(n2485), .A2(n2333), .ZN(n2487) );
  NAND2_X1 U469 ( .A1(n2485), .A2(n2343), .ZN(n2496) );
  NAND2_X1 U470 ( .A1(n2485), .A2(n2353), .ZN(n2505) );
  NAND2_X1 U471 ( .A1(n2485), .A2(n2363), .ZN(n2514) );
  NAND2_X1 U472 ( .A1(n2485), .A2(n2373), .ZN(n2523) );
  NAND2_X1 U473 ( .A1(n2485), .A2(n2383), .ZN(n2532) );
  NAND2_X1 U474 ( .A1(n2485), .A2(n2393), .ZN(n2541) );
  NAND2_X1 U475 ( .A1(n2485), .A2(n2403), .ZN(n2550) );
  NAND2_X1 U476 ( .A1(n2485), .A2(n2413), .ZN(n2559) );
  NAND2_X1 U477 ( .A1(n2485), .A2(n2423), .ZN(n2568) );
  NAND2_X1 U478 ( .A1(n2485), .A2(n2433), .ZN(n2577) );
  NAND2_X1 U479 ( .A1(n2485), .A2(n2443), .ZN(n2586) );
  NAND2_X1 U480 ( .A1(n2485), .A2(n2453), .ZN(n2595) );
  NAND2_X1 U481 ( .A1(n2485), .A2(n2463), .ZN(n2604) );
  NAND2_X1 U482 ( .A1(n2485), .A2(n2473), .ZN(n2613) );
  NAND2_X1 U483 ( .A1(n2631), .A2(n2322), .ZN(n2623) );
  NAND2_X1 U484 ( .A1(n2631), .A2(n2333), .ZN(n2633) );
  NAND2_X1 U485 ( .A1(n2631), .A2(n2343), .ZN(n2642) );
  NAND2_X1 U486 ( .A1(n2631), .A2(n2353), .ZN(n2651) );
  NAND2_X1 U487 ( .A1(n2631), .A2(n2363), .ZN(n2660) );
  NAND2_X1 U488 ( .A1(n2631), .A2(n2373), .ZN(n2669) );
  NAND2_X1 U489 ( .A1(n2631), .A2(n2383), .ZN(n2678) );
  NAND2_X1 U490 ( .A1(n2631), .A2(n2393), .ZN(n2687) );
  NAND2_X1 U491 ( .A1(n2631), .A2(n2403), .ZN(n2696) );
  NAND2_X1 U492 ( .A1(n2631), .A2(n2413), .ZN(n2705) );
  NAND2_X1 U493 ( .A1(n2631), .A2(n2423), .ZN(n2714) );
  NAND2_X1 U494 ( .A1(n2631), .A2(n2433), .ZN(n2723) );
  NAND2_X1 U495 ( .A1(n2631), .A2(n2443), .ZN(n2732) );
  NAND2_X1 U496 ( .A1(n2631), .A2(n2453), .ZN(n2741) );
  NAND2_X1 U497 ( .A1(n2631), .A2(n2463), .ZN(n2750) );
  NAND2_X1 U498 ( .A1(n2631), .A2(n2473), .ZN(n2759) );
  NAND2_X1 U499 ( .A1(n2777), .A2(n2322), .ZN(n2769) );
  NAND2_X1 U500 ( .A1(n2777), .A2(n2333), .ZN(n2779) );
  NAND2_X1 U501 ( .A1(n2777), .A2(n2343), .ZN(n2788) );
  NAND2_X1 U502 ( .A1(n2777), .A2(n2353), .ZN(n2797) );
  NAND2_X1 U503 ( .A1(n2777), .A2(n2363), .ZN(n2806) );
  NAND2_X1 U504 ( .A1(n2777), .A2(n2373), .ZN(n2815) );
  NAND2_X1 U505 ( .A1(n2777), .A2(n2383), .ZN(n2824) );
  NAND2_X1 U506 ( .A1(n2777), .A2(n2393), .ZN(n2833) );
  NAND2_X1 U507 ( .A1(n2777), .A2(n2403), .ZN(n2842) );
  NAND2_X1 U508 ( .A1(n2777), .A2(n2413), .ZN(n2851) );
  NAND2_X1 U509 ( .A1(n2777), .A2(n2423), .ZN(n2860) );
  NAND2_X1 U510 ( .A1(n2777), .A2(n2433), .ZN(n2869) );
  NAND2_X1 U511 ( .A1(n2777), .A2(n2443), .ZN(n2878) );
  NAND2_X1 U512 ( .A1(n2777), .A2(n2453), .ZN(n2887) );
  NAND2_X1 U513 ( .A1(n2777), .A2(n2463), .ZN(n2896) );
  NAND2_X1 U514 ( .A1(n2777), .A2(n2473), .ZN(n2905) );
  NAND2_X1 U515 ( .A1(n4085), .A2(n2322), .ZN(n4077) );
  NAND2_X1 U516 ( .A1(n4085), .A2(n2333), .ZN(n4087) );
  NAND2_X1 U517 ( .A1(n4085), .A2(n2343), .ZN(n4096) );
  NAND2_X1 U518 ( .A1(n4085), .A2(n2353), .ZN(n4105) );
  NAND2_X1 U519 ( .A1(n4085), .A2(n2363), .ZN(n4114) );
  NAND2_X1 U520 ( .A1(n4085), .A2(n2373), .ZN(n4123) );
  NAND2_X1 U521 ( .A1(n4085), .A2(n2383), .ZN(n4132) );
  NAND2_X1 U522 ( .A1(n4085), .A2(n2393), .ZN(n4141) );
  NAND2_X1 U523 ( .A1(n4085), .A2(n2403), .ZN(n4150) );
  NAND2_X1 U524 ( .A1(n4085), .A2(n2413), .ZN(n4159) );
  NAND2_X1 U525 ( .A1(n4085), .A2(n2423), .ZN(n4168) );
  NAND2_X1 U526 ( .A1(n4085), .A2(n2433), .ZN(n4177) );
  NAND2_X1 U527 ( .A1(n4085), .A2(n2443), .ZN(n4186) );
  NAND2_X1 U528 ( .A1(n4085), .A2(n2453), .ZN(n4195) );
  NAND2_X1 U529 ( .A1(n4085), .A2(n2463), .ZN(n4204) );
  NAND2_X1 U530 ( .A1(n4085), .A2(n2473), .ZN(n4213) );
  BUF_X1 U531 ( .A(addr_r[0]), .Z(n6743) );
  BUF_X1 U532 ( .A(n6741), .Z(n6744) );
  BUF_X1 U533 ( .A(addr_r[0]), .Z(n6745) );
  BUF_X1 U534 ( .A(n6742), .Z(n6752) );
  BUF_X1 U535 ( .A(n6742), .Z(n6755) );
  BUF_X1 U536 ( .A(n6742), .Z(n6753) );
  BUF_X1 U537 ( .A(n6742), .Z(n6754) );
  BUF_X1 U538 ( .A(n6741), .Z(n6763) );
  BUF_X1 U539 ( .A(n6741), .Z(n6764) );
  BUF_X1 U540 ( .A(n6741), .Z(n6765) );
  BUF_X1 U541 ( .A(n6741), .Z(n6766) );
  BUF_X1 U542 ( .A(n6740), .Z(n6774) );
  BUF_X1 U543 ( .A(n6740), .Z(n6775) );
  BUF_X1 U544 ( .A(n6740), .Z(n6776) );
  BUF_X1 U545 ( .A(n6740), .Z(n6777) );
  BUF_X1 U546 ( .A(n6721), .Z(n6722) );
  BUF_X1 U547 ( .A(n6721), .Z(n6723) );
  BUF_X1 U548 ( .A(n6721), .Z(n6724) );
  BUF_X1 U549 ( .A(n6721), .Z(n6725) );
  BUF_X1 U550 ( .A(n6720), .Z(n6726) );
  BUF_X1 U551 ( .A(n6720), .Z(n6727) );
  BUF_X1 U552 ( .A(n6720), .Z(n6728) );
  BUF_X1 U553 ( .A(n6720), .Z(n6729) );
  BUF_X1 U554 ( .A(n6720), .Z(n6730) );
  BUF_X1 U555 ( .A(n6719), .Z(n6731) );
  BUF_X1 U556 ( .A(n6719), .Z(n6732) );
  BUF_X1 U557 ( .A(n6719), .Z(n6733) );
  BUF_X1 U558 ( .A(n6719), .Z(n6734) );
  BUF_X1 U559 ( .A(n6719), .Z(n6735) );
  BUF_X1 U560 ( .A(n6718), .Z(n6738) );
  BUF_X1 U561 ( .A(n6718), .Z(n6737) );
  BUF_X1 U562 ( .A(n6718), .Z(n6736) );
  AND3_X1 U563 ( .A1(we_s), .A2(n2475), .A3(n3059), .ZN(n2923) );
  AND3_X1 U564 ( .A1(n2621), .A2(we_s), .A3(n3059), .ZN(n3069) );
  AND3_X1 U565 ( .A1(n2767), .A2(we_s), .A3(n3059), .ZN(n3214) );
  AND3_X1 U566 ( .A1(n2913), .A2(we_s), .A3(n3059), .ZN(n3359) );
  AND3_X1 U567 ( .A1(we_s), .A2(n2475), .A3(n3640), .ZN(n3504) );
  AND3_X1 U568 ( .A1(n2621), .A2(we_s), .A3(n3640), .ZN(n3650) );
  AND3_X1 U569 ( .A1(n2767), .A2(we_s), .A3(n3640), .ZN(n3795) );
  AND3_X1 U570 ( .A1(n2913), .A2(we_s), .A3(n3640), .ZN(n3940) );
  AND3_X1 U571 ( .A1(n2621), .A2(we_s), .A3(n4221), .ZN(n4231) );
  AND3_X1 U572 ( .A1(n2767), .A2(we_s), .A3(n4221), .ZN(n4376) );
  AND3_X1 U573 ( .A1(n2913), .A2(we_s), .A3(n4221), .ZN(n4521) );
  AND3_X1 U574 ( .A1(we_s), .A2(n2474), .A3(n2621), .ZN(n2485) );
  AND3_X1 U575 ( .A1(we_s), .A2(n2474), .A3(n2767), .ZN(n2631) );
  AND3_X1 U576 ( .A1(we_s), .A2(n2474), .A3(n2913), .ZN(n2777) );
  AND3_X1 U577 ( .A1(we_s), .A2(n2475), .A3(n4221), .ZN(n4085) );
  NOR2_X1 U578 ( .A1(n9089), .A2(n7936), .ZN(n4523) );
  NOR2_X1 U579 ( .A1(n9091), .A2(n9090), .ZN(n4522) );
  NOR2_X1 U580 ( .A1(n9095), .A2(n9094), .ZN(n2474) );
  BUF_X1 U581 ( .A(n6717), .Z(n6707) );
  BUF_X1 U582 ( .A(n6717), .Z(n6708) );
  BUF_X1 U583 ( .A(n6717), .Z(n6709) );
  BUF_X1 U584 ( .A(n6717), .Z(n6710) );
  BUF_X1 U585 ( .A(n6700), .Z(n6698) );
  BUF_X1 U586 ( .A(addr_r[4]), .Z(n6699) );
  NOR2_X1 U587 ( .A1(n9093), .A2(n9092), .ZN(n2475) );
  BUF_X1 U588 ( .A(n6739), .Z(n6718) );
  BUF_X1 U589 ( .A(addr_r[1]), .Z(n6721) );
  BUF_X1 U590 ( .A(n6739), .Z(n6720) );
  BUF_X1 U591 ( .A(n6739), .Z(n6719) );
  BUF_X1 U592 ( .A(addr_r[0]), .Z(n6742) );
  BUF_X1 U593 ( .A(n6783), .Z(n6741) );
  BUF_X1 U594 ( .A(n6783), .Z(n6740) );
  NOR2_X1 U595 ( .A1(addr_w[0]), .A2(addr_w[1]), .ZN(n4553) );
  NOR2_X1 U596 ( .A1(n7936), .A2(addr_w[1]), .ZN(n4543) );
  NOR2_X1 U597 ( .A1(n9089), .A2(addr_w[0]), .ZN(n4533) );
  NOR2_X1 U598 ( .A1(addr_w[2]), .A2(addr_w[3]), .ZN(n4637) );
  NOR2_X1 U599 ( .A1(n9091), .A2(addr_w[2]), .ZN(n4563) );
  NOR2_X1 U600 ( .A1(n9090), .A2(addr_w[3]), .ZN(n4600) );
  BUF_X1 U601 ( .A(addr_r[3]), .Z(n6701) );
  BUF_X1 U602 ( .A(addr_r[5]), .Z(n6697) );
  NOR2_X1 U603 ( .A1(addr_w[6]), .A2(addr_w[7]), .ZN(n4221) );
  NOR2_X1 U604 ( .A1(addr_w[4]), .A2(addr_w[5]), .ZN(n2913) );
  NOR2_X1 U605 ( .A1(n9092), .A2(addr_w[5]), .ZN(n2767) );
  NOR2_X1 U606 ( .A1(n9093), .A2(addr_w[4]), .ZN(n2621) );
  NOR2_X1 U607 ( .A1(n9095), .A2(addr_w[6]), .ZN(n3059) );
  NOR2_X1 U608 ( .A1(n9094), .A2(addr_w[7]), .ZN(n3640) );
  INV_X1 U609 ( .A(addr_w[1]), .ZN(n9089) );
  INV_X1 U610 ( .A(addr_w[0]), .ZN(n7936) );
  INV_X1 U611 ( .A(addr_w[2]), .ZN(n9090) );
  INV_X1 U612 ( .A(addr_w[3]), .ZN(n9091) );
  INV_X1 U613 ( .A(addr_w[6]), .ZN(n9094) );
  INV_X1 U614 ( .A(addr_w[4]), .ZN(n9092) );
  INV_X1 U615 ( .A(addr_w[5]), .ZN(n9093) );
  BUF_X1 U616 ( .A(addr_r[2]), .Z(n6717) );
  INV_X1 U617 ( .A(addr_w[7]), .ZN(n9095) );
  BUF_X1 U618 ( .A(addr_r[1]), .Z(n6739) );
  BUF_X1 U619 ( .A(addr_r[0]), .Z(n6783) );
  INV_X1 U620 ( .A(n3459), .ZN(n6856) );
  AOI22_X1 U621 ( .A1(reg_mem[992]), .A2(n3460), .B1(n6864), .B2(data_w[0]), 
        .ZN(n3459) );
  INV_X1 U622 ( .A(n3461), .ZN(n6857) );
  AOI22_X1 U623 ( .A1(reg_mem[993]), .A2(n3460), .B1(n6864), .B2(data_w[1]), 
        .ZN(n3461) );
  INV_X1 U624 ( .A(n3462), .ZN(n6858) );
  AOI22_X1 U625 ( .A1(reg_mem[994]), .A2(n3460), .B1(n6864), .B2(data_w[2]), 
        .ZN(n3462) );
  INV_X1 U626 ( .A(n3463), .ZN(n6859) );
  AOI22_X1 U627 ( .A1(reg_mem[995]), .A2(n3460), .B1(n6864), .B2(data_w[3]), 
        .ZN(n3463) );
  INV_X1 U628 ( .A(n3464), .ZN(n6860) );
  AOI22_X1 U629 ( .A1(reg_mem[996]), .A2(n3460), .B1(n6864), .B2(data_w[4]), 
        .ZN(n3464) );
  INV_X1 U630 ( .A(n3465), .ZN(n6861) );
  AOI22_X1 U631 ( .A1(reg_mem[997]), .A2(n3460), .B1(n6864), .B2(data_w[5]), 
        .ZN(n3465) );
  INV_X1 U632 ( .A(n3466), .ZN(n6862) );
  AOI22_X1 U633 ( .A1(reg_mem[998]), .A2(n3460), .B1(n6864), .B2(data_w[6]), 
        .ZN(n3466) );
  INV_X1 U634 ( .A(n3467), .ZN(n6863) );
  AOI22_X1 U635 ( .A1(reg_mem[999]), .A2(n3460), .B1(n6864), .B2(data_w[7]), 
        .ZN(n3467) );
  INV_X1 U636 ( .A(n3468), .ZN(n8585) );
  AOI22_X1 U637 ( .A1(reg_mem[1000]), .A2(n3469), .B1(n8593), .B2(data_w[0]), 
        .ZN(n3468) );
  INV_X1 U638 ( .A(n3470), .ZN(n8586) );
  AOI22_X1 U639 ( .A1(reg_mem[1001]), .A2(n3469), .B1(n8593), .B2(data_w[1]), 
        .ZN(n3470) );
  INV_X1 U640 ( .A(n3471), .ZN(n8587) );
  AOI22_X1 U641 ( .A1(reg_mem[1002]), .A2(n3469), .B1(n8593), .B2(data_w[2]), 
        .ZN(n3471) );
  INV_X1 U642 ( .A(n3472), .ZN(n8588) );
  AOI22_X1 U643 ( .A1(reg_mem[1003]), .A2(n3469), .B1(n8593), .B2(data_w[3]), 
        .ZN(n3472) );
  INV_X1 U644 ( .A(n3473), .ZN(n8589) );
  AOI22_X1 U645 ( .A1(reg_mem[1004]), .A2(n3469), .B1(n8593), .B2(data_w[4]), 
        .ZN(n3473) );
  INV_X1 U646 ( .A(n3474), .ZN(n8590) );
  AOI22_X1 U647 ( .A1(reg_mem[1005]), .A2(n3469), .B1(n8593), .B2(data_w[5]), 
        .ZN(n3474) );
  INV_X1 U648 ( .A(n3475), .ZN(n8591) );
  AOI22_X1 U649 ( .A1(reg_mem[1006]), .A2(n3469), .B1(n8593), .B2(data_w[6]), 
        .ZN(n3475) );
  INV_X1 U650 ( .A(n3476), .ZN(n8592) );
  AOI22_X1 U651 ( .A1(reg_mem[1007]), .A2(n3469), .B1(n8593), .B2(data_w[7]), 
        .ZN(n3476) );
  INV_X1 U652 ( .A(n3477), .ZN(n7432) );
  AOI22_X1 U653 ( .A1(reg_mem[1008]), .A2(n3478), .B1(n7440), .B2(data_w[0]), 
        .ZN(n3477) );
  INV_X1 U654 ( .A(n3479), .ZN(n7433) );
  AOI22_X1 U655 ( .A1(reg_mem[1009]), .A2(n3478), .B1(n7440), .B2(data_w[1]), 
        .ZN(n3479) );
  INV_X1 U656 ( .A(n3480), .ZN(n7434) );
  AOI22_X1 U657 ( .A1(reg_mem[1010]), .A2(n3478), .B1(n7440), .B2(data_w[2]), 
        .ZN(n3480) );
  INV_X1 U658 ( .A(n3481), .ZN(n7435) );
  AOI22_X1 U659 ( .A1(reg_mem[1011]), .A2(n3478), .B1(n7440), .B2(data_w[3]), 
        .ZN(n3481) );
  INV_X1 U660 ( .A(n3482), .ZN(n7436) );
  AOI22_X1 U661 ( .A1(reg_mem[1012]), .A2(n3478), .B1(n7440), .B2(data_w[4]), 
        .ZN(n3482) );
  INV_X1 U662 ( .A(n3483), .ZN(n7437) );
  AOI22_X1 U663 ( .A1(reg_mem[1013]), .A2(n3478), .B1(n7440), .B2(data_w[5]), 
        .ZN(n3483) );
  INV_X1 U664 ( .A(n3484), .ZN(n7438) );
  AOI22_X1 U665 ( .A1(reg_mem[1014]), .A2(n3478), .B1(n7440), .B2(data_w[6]), 
        .ZN(n3484) );
  INV_X1 U666 ( .A(n3485), .ZN(n7439) );
  AOI22_X1 U667 ( .A1(reg_mem[1015]), .A2(n3478), .B1(n7440), .B2(data_w[7]), 
        .ZN(n3485) );
  INV_X1 U668 ( .A(n3486), .ZN(n8009) );
  AOI22_X1 U669 ( .A1(reg_mem[1016]), .A2(n3487), .B1(n8017), .B2(data_w[0]), 
        .ZN(n3486) );
  INV_X1 U670 ( .A(n3488), .ZN(n8010) );
  AOI22_X1 U671 ( .A1(reg_mem[1017]), .A2(n3487), .B1(n8017), .B2(data_w[1]), 
        .ZN(n3488) );
  INV_X1 U672 ( .A(n3489), .ZN(n8011) );
  AOI22_X1 U673 ( .A1(reg_mem[1018]), .A2(n3487), .B1(n8017), .B2(data_w[2]), 
        .ZN(n3489) );
  INV_X1 U674 ( .A(n3490), .ZN(n8012) );
  AOI22_X1 U675 ( .A1(reg_mem[1019]), .A2(n3487), .B1(n8017), .B2(data_w[3]), 
        .ZN(n3490) );
  INV_X1 U676 ( .A(n3491), .ZN(n8013) );
  AOI22_X1 U677 ( .A1(reg_mem[1020]), .A2(n3487), .B1(n8017), .B2(data_w[4]), 
        .ZN(n3491) );
  INV_X1 U678 ( .A(n3492), .ZN(n8014) );
  AOI22_X1 U679 ( .A1(reg_mem[1021]), .A2(n3487), .B1(n8017), .B2(data_w[5]), 
        .ZN(n3492) );
  INV_X1 U680 ( .A(n3493), .ZN(n8015) );
  AOI22_X1 U681 ( .A1(reg_mem[1022]), .A2(n3487), .B1(n8017), .B2(data_w[6]), 
        .ZN(n3493) );
  INV_X1 U682 ( .A(n3494), .ZN(n8016) );
  AOI22_X1 U683 ( .A1(reg_mem[1023]), .A2(n3487), .B1(n8017), .B2(data_w[7]), 
        .ZN(n3494) );
  INV_X1 U684 ( .A(n3495), .ZN(n7279) );
  AOI22_X1 U685 ( .A1(reg_mem[1024]), .A2(n3496), .B1(n7287), .B2(data_w[0]), 
        .ZN(n3495) );
  INV_X1 U686 ( .A(n3497), .ZN(n7280) );
  AOI22_X1 U687 ( .A1(reg_mem[1025]), .A2(n3496), .B1(n7287), .B2(data_w[1]), 
        .ZN(n3497) );
  INV_X1 U688 ( .A(n3498), .ZN(n7281) );
  AOI22_X1 U689 ( .A1(reg_mem[1026]), .A2(n3496), .B1(n7287), .B2(data_w[2]), 
        .ZN(n3498) );
  INV_X1 U690 ( .A(n3499), .ZN(n7282) );
  AOI22_X1 U691 ( .A1(reg_mem[1027]), .A2(n3496), .B1(n7287), .B2(data_w[3]), 
        .ZN(n3499) );
  INV_X1 U692 ( .A(n3500), .ZN(n7283) );
  AOI22_X1 U693 ( .A1(reg_mem[1028]), .A2(n3496), .B1(n7287), .B2(data_w[4]), 
        .ZN(n3500) );
  INV_X1 U694 ( .A(n3501), .ZN(n7284) );
  AOI22_X1 U695 ( .A1(reg_mem[1029]), .A2(n3496), .B1(n7287), .B2(data_w[5]), 
        .ZN(n3501) );
  INV_X1 U696 ( .A(n3502), .ZN(n7285) );
  AOI22_X1 U697 ( .A1(reg_mem[1030]), .A2(n3496), .B1(n7287), .B2(data_w[6]), 
        .ZN(n3502) );
  INV_X1 U698 ( .A(n3503), .ZN(n7286) );
  AOI22_X1 U699 ( .A1(reg_mem[1031]), .A2(n3496), .B1(n7287), .B2(data_w[7]), 
        .ZN(n3503) );
  INV_X1 U700 ( .A(n3505), .ZN(n9008) );
  AOI22_X1 U701 ( .A1(reg_mem[1032]), .A2(n3506), .B1(n9016), .B2(data_w[0]), 
        .ZN(n3505) );
  INV_X1 U702 ( .A(n3507), .ZN(n9009) );
  AOI22_X1 U703 ( .A1(reg_mem[1033]), .A2(n3506), .B1(n9016), .B2(data_w[1]), 
        .ZN(n3507) );
  INV_X1 U704 ( .A(n3508), .ZN(n9010) );
  AOI22_X1 U705 ( .A1(reg_mem[1034]), .A2(n3506), .B1(n9016), .B2(data_w[2]), 
        .ZN(n3508) );
  INV_X1 U706 ( .A(n3509), .ZN(n9011) );
  AOI22_X1 U707 ( .A1(reg_mem[1035]), .A2(n3506), .B1(n9016), .B2(data_w[3]), 
        .ZN(n3509) );
  INV_X1 U708 ( .A(n3510), .ZN(n9012) );
  AOI22_X1 U709 ( .A1(reg_mem[1036]), .A2(n3506), .B1(n9016), .B2(data_w[4]), 
        .ZN(n3510) );
  INV_X1 U710 ( .A(n3511), .ZN(n9013) );
  AOI22_X1 U711 ( .A1(reg_mem[1037]), .A2(n3506), .B1(n9016), .B2(data_w[5]), 
        .ZN(n3511) );
  INV_X1 U712 ( .A(n3512), .ZN(n9014) );
  AOI22_X1 U713 ( .A1(reg_mem[1038]), .A2(n3506), .B1(n9016), .B2(data_w[6]), 
        .ZN(n3512) );
  INV_X1 U714 ( .A(n3513), .ZN(n9015) );
  AOI22_X1 U715 ( .A1(reg_mem[1039]), .A2(n3506), .B1(n9016), .B2(data_w[7]), 
        .ZN(n3513) );
  INV_X1 U716 ( .A(n3514), .ZN(n7855) );
  AOI22_X1 U717 ( .A1(reg_mem[1040]), .A2(n3515), .B1(n7863), .B2(data_w[0]), 
        .ZN(n3514) );
  INV_X1 U718 ( .A(n3516), .ZN(n7856) );
  AOI22_X1 U719 ( .A1(reg_mem[1041]), .A2(n3515), .B1(n7863), .B2(data_w[1]), 
        .ZN(n3516) );
  INV_X1 U720 ( .A(n3517), .ZN(n7857) );
  AOI22_X1 U721 ( .A1(reg_mem[1042]), .A2(n3515), .B1(n7863), .B2(data_w[2]), 
        .ZN(n3517) );
  INV_X1 U722 ( .A(n3518), .ZN(n7858) );
  AOI22_X1 U723 ( .A1(reg_mem[1043]), .A2(n3515), .B1(n7863), .B2(data_w[3]), 
        .ZN(n3518) );
  INV_X1 U724 ( .A(n3519), .ZN(n7859) );
  AOI22_X1 U725 ( .A1(reg_mem[1044]), .A2(n3515), .B1(n7863), .B2(data_w[4]), 
        .ZN(n3519) );
  INV_X1 U726 ( .A(n3520), .ZN(n7860) );
  AOI22_X1 U727 ( .A1(reg_mem[1045]), .A2(n3515), .B1(n7863), .B2(data_w[5]), 
        .ZN(n3520) );
  INV_X1 U728 ( .A(n3521), .ZN(n7861) );
  AOI22_X1 U729 ( .A1(reg_mem[1046]), .A2(n3515), .B1(n7863), .B2(data_w[6]), 
        .ZN(n3521) );
  INV_X1 U730 ( .A(n3522), .ZN(n7862) );
  AOI22_X1 U731 ( .A1(reg_mem[1047]), .A2(n3515), .B1(n7863), .B2(data_w[7]), 
        .ZN(n3522) );
  INV_X1 U732 ( .A(n3523), .ZN(n8432) );
  AOI22_X1 U733 ( .A1(reg_mem[1048]), .A2(n3524), .B1(n8440), .B2(data_w[0]), 
        .ZN(n3523) );
  INV_X1 U734 ( .A(n3525), .ZN(n8433) );
  AOI22_X1 U735 ( .A1(reg_mem[1049]), .A2(n3524), .B1(n8440), .B2(data_w[1]), 
        .ZN(n3525) );
  INV_X1 U736 ( .A(n3526), .ZN(n8434) );
  AOI22_X1 U737 ( .A1(reg_mem[1050]), .A2(n3524), .B1(n8440), .B2(data_w[2]), 
        .ZN(n3526) );
  INV_X1 U738 ( .A(n3527), .ZN(n8435) );
  AOI22_X1 U739 ( .A1(reg_mem[1051]), .A2(n3524), .B1(n8440), .B2(data_w[3]), 
        .ZN(n3527) );
  INV_X1 U740 ( .A(n3528), .ZN(n8436) );
  AOI22_X1 U741 ( .A1(reg_mem[1052]), .A2(n3524), .B1(n8440), .B2(data_w[4]), 
        .ZN(n3528) );
  INV_X1 U742 ( .A(n3529), .ZN(n8437) );
  AOI22_X1 U743 ( .A1(reg_mem[1053]), .A2(n3524), .B1(n8440), .B2(data_w[5]), 
        .ZN(n3529) );
  INV_X1 U744 ( .A(n3530), .ZN(n8438) );
  AOI22_X1 U745 ( .A1(reg_mem[1054]), .A2(n3524), .B1(n8440), .B2(data_w[6]), 
        .ZN(n3530) );
  INV_X1 U746 ( .A(n3531), .ZN(n8439) );
  AOI22_X1 U747 ( .A1(reg_mem[1055]), .A2(n3524), .B1(n8440), .B2(data_w[7]), 
        .ZN(n3531) );
  INV_X1 U748 ( .A(n3532), .ZN(n7135) );
  AOI22_X1 U749 ( .A1(reg_mem[1056]), .A2(n3533), .B1(n7143), .B2(data_w[0]), 
        .ZN(n3532) );
  INV_X1 U750 ( .A(n3534), .ZN(n7136) );
  AOI22_X1 U751 ( .A1(reg_mem[1057]), .A2(n3533), .B1(n7143), .B2(data_w[1]), 
        .ZN(n3534) );
  INV_X1 U752 ( .A(n3535), .ZN(n7137) );
  AOI22_X1 U753 ( .A1(reg_mem[1058]), .A2(n3533), .B1(n7143), .B2(data_w[2]), 
        .ZN(n3535) );
  INV_X1 U754 ( .A(n3536), .ZN(n7138) );
  AOI22_X1 U755 ( .A1(reg_mem[1059]), .A2(n3533), .B1(n7143), .B2(data_w[3]), 
        .ZN(n3536) );
  INV_X1 U756 ( .A(n3537), .ZN(n7139) );
  AOI22_X1 U757 ( .A1(reg_mem[1060]), .A2(n3533), .B1(n7143), .B2(data_w[4]), 
        .ZN(n3537) );
  INV_X1 U758 ( .A(n3538), .ZN(n7140) );
  AOI22_X1 U759 ( .A1(reg_mem[1061]), .A2(n3533), .B1(n7143), .B2(data_w[5]), 
        .ZN(n3538) );
  INV_X1 U760 ( .A(n3539), .ZN(n7141) );
  AOI22_X1 U761 ( .A1(reg_mem[1062]), .A2(n3533), .B1(n7143), .B2(data_w[6]), 
        .ZN(n3539) );
  INV_X1 U762 ( .A(n3540), .ZN(n7142) );
  AOI22_X1 U763 ( .A1(reg_mem[1063]), .A2(n3533), .B1(n7143), .B2(data_w[7]), 
        .ZN(n3540) );
  INV_X1 U764 ( .A(n3541), .ZN(n8864) );
  AOI22_X1 U765 ( .A1(reg_mem[1064]), .A2(n3542), .B1(n8872), .B2(data_w[0]), 
        .ZN(n3541) );
  INV_X1 U766 ( .A(n3543), .ZN(n8865) );
  AOI22_X1 U767 ( .A1(reg_mem[1065]), .A2(n3542), .B1(n8872), .B2(data_w[1]), 
        .ZN(n3543) );
  INV_X1 U768 ( .A(n3544), .ZN(n8866) );
  AOI22_X1 U769 ( .A1(reg_mem[1066]), .A2(n3542), .B1(n8872), .B2(data_w[2]), 
        .ZN(n3544) );
  INV_X1 U770 ( .A(n3545), .ZN(n8867) );
  AOI22_X1 U771 ( .A1(reg_mem[1067]), .A2(n3542), .B1(n8872), .B2(data_w[3]), 
        .ZN(n3545) );
  INV_X1 U772 ( .A(n3546), .ZN(n8868) );
  AOI22_X1 U773 ( .A1(reg_mem[1068]), .A2(n3542), .B1(n8872), .B2(data_w[4]), 
        .ZN(n3546) );
  INV_X1 U774 ( .A(n3547), .ZN(n8869) );
  AOI22_X1 U775 ( .A1(reg_mem[1069]), .A2(n3542), .B1(n8872), .B2(data_w[5]), 
        .ZN(n3547) );
  INV_X1 U776 ( .A(n3548), .ZN(n8870) );
  AOI22_X1 U777 ( .A1(reg_mem[1070]), .A2(n3542), .B1(n8872), .B2(data_w[6]), 
        .ZN(n3548) );
  INV_X1 U778 ( .A(n3549), .ZN(n8871) );
  AOI22_X1 U779 ( .A1(reg_mem[1071]), .A2(n3542), .B1(n8872), .B2(data_w[7]), 
        .ZN(n3549) );
  INV_X1 U780 ( .A(n3550), .ZN(n7711) );
  AOI22_X1 U781 ( .A1(reg_mem[1072]), .A2(n3551), .B1(n7719), .B2(data_w[0]), 
        .ZN(n3550) );
  INV_X1 U782 ( .A(n3552), .ZN(n7712) );
  AOI22_X1 U783 ( .A1(reg_mem[1073]), .A2(n3551), .B1(n7719), .B2(data_w[1]), 
        .ZN(n3552) );
  INV_X1 U784 ( .A(n3553), .ZN(n7713) );
  AOI22_X1 U785 ( .A1(reg_mem[1074]), .A2(n3551), .B1(n7719), .B2(data_w[2]), 
        .ZN(n3553) );
  INV_X1 U786 ( .A(n3554), .ZN(n7714) );
  AOI22_X1 U787 ( .A1(reg_mem[1075]), .A2(n3551), .B1(n7719), .B2(data_w[3]), 
        .ZN(n3554) );
  INV_X1 U788 ( .A(n3555), .ZN(n7715) );
  AOI22_X1 U789 ( .A1(reg_mem[1076]), .A2(n3551), .B1(n7719), .B2(data_w[4]), 
        .ZN(n3555) );
  INV_X1 U790 ( .A(n3556), .ZN(n7716) );
  AOI22_X1 U791 ( .A1(reg_mem[1077]), .A2(n3551), .B1(n7719), .B2(data_w[5]), 
        .ZN(n3556) );
  INV_X1 U792 ( .A(n3557), .ZN(n7717) );
  AOI22_X1 U793 ( .A1(reg_mem[1078]), .A2(n3551), .B1(n7719), .B2(data_w[6]), 
        .ZN(n3557) );
  INV_X1 U794 ( .A(n3558), .ZN(n7718) );
  AOI22_X1 U795 ( .A1(reg_mem[1079]), .A2(n3551), .B1(n7719), .B2(data_w[7]), 
        .ZN(n3558) );
  INV_X1 U796 ( .A(n3559), .ZN(n8288) );
  AOI22_X1 U797 ( .A1(reg_mem[1080]), .A2(n3560), .B1(n8296), .B2(data_w[0]), 
        .ZN(n3559) );
  INV_X1 U798 ( .A(n3561), .ZN(n8289) );
  AOI22_X1 U799 ( .A1(reg_mem[1081]), .A2(n3560), .B1(n8296), .B2(data_w[1]), 
        .ZN(n3561) );
  INV_X1 U800 ( .A(n3562), .ZN(n8290) );
  AOI22_X1 U801 ( .A1(reg_mem[1082]), .A2(n3560), .B1(n8296), .B2(data_w[2]), 
        .ZN(n3562) );
  INV_X1 U802 ( .A(n3563), .ZN(n8291) );
  AOI22_X1 U803 ( .A1(reg_mem[1083]), .A2(n3560), .B1(n8296), .B2(data_w[3]), 
        .ZN(n3563) );
  INV_X1 U804 ( .A(n3564), .ZN(n8292) );
  AOI22_X1 U805 ( .A1(reg_mem[1084]), .A2(n3560), .B1(n8296), .B2(data_w[4]), 
        .ZN(n3564) );
  INV_X1 U806 ( .A(n3565), .ZN(n8293) );
  AOI22_X1 U807 ( .A1(reg_mem[1085]), .A2(n3560), .B1(n8296), .B2(data_w[5]), 
        .ZN(n3565) );
  INV_X1 U808 ( .A(n3566), .ZN(n8294) );
  AOI22_X1 U809 ( .A1(reg_mem[1086]), .A2(n3560), .B1(n8296), .B2(data_w[6]), 
        .ZN(n3566) );
  INV_X1 U810 ( .A(n3567), .ZN(n8295) );
  AOI22_X1 U811 ( .A1(reg_mem[1087]), .A2(n3560), .B1(n8296), .B2(data_w[7]), 
        .ZN(n3567) );
  INV_X1 U812 ( .A(n3568), .ZN(n6991) );
  AOI22_X1 U813 ( .A1(reg_mem[1088]), .A2(n3569), .B1(n6999), .B2(data_w[0]), 
        .ZN(n3568) );
  INV_X1 U814 ( .A(n3570), .ZN(n6992) );
  AOI22_X1 U815 ( .A1(reg_mem[1089]), .A2(n3569), .B1(n6999), .B2(data_w[1]), 
        .ZN(n3570) );
  INV_X1 U816 ( .A(n3571), .ZN(n6993) );
  AOI22_X1 U817 ( .A1(reg_mem[1090]), .A2(n3569), .B1(n6999), .B2(data_w[2]), 
        .ZN(n3571) );
  INV_X1 U818 ( .A(n3572), .ZN(n6994) );
  AOI22_X1 U819 ( .A1(reg_mem[1091]), .A2(n3569), .B1(n6999), .B2(data_w[3]), 
        .ZN(n3572) );
  INV_X1 U820 ( .A(n3573), .ZN(n6995) );
  AOI22_X1 U821 ( .A1(reg_mem[1092]), .A2(n3569), .B1(n6999), .B2(data_w[4]), 
        .ZN(n3573) );
  INV_X1 U822 ( .A(n3574), .ZN(n6996) );
  AOI22_X1 U823 ( .A1(reg_mem[1093]), .A2(n3569), .B1(n6999), .B2(data_w[5]), 
        .ZN(n3574) );
  INV_X1 U824 ( .A(n3575), .ZN(n6997) );
  AOI22_X1 U825 ( .A1(reg_mem[1094]), .A2(n3569), .B1(n6999), .B2(data_w[6]), 
        .ZN(n3575) );
  INV_X1 U826 ( .A(n3576), .ZN(n6998) );
  AOI22_X1 U827 ( .A1(reg_mem[1095]), .A2(n3569), .B1(n6999), .B2(data_w[7]), 
        .ZN(n3576) );
  INV_X1 U828 ( .A(n3577), .ZN(n8720) );
  AOI22_X1 U829 ( .A1(reg_mem[1096]), .A2(n3578), .B1(n8728), .B2(data_w[0]), 
        .ZN(n3577) );
  INV_X1 U830 ( .A(n3579), .ZN(n8721) );
  AOI22_X1 U831 ( .A1(reg_mem[1097]), .A2(n3578), .B1(n8728), .B2(data_w[1]), 
        .ZN(n3579) );
  INV_X1 U832 ( .A(n3580), .ZN(n8722) );
  AOI22_X1 U833 ( .A1(reg_mem[1098]), .A2(n3578), .B1(n8728), .B2(data_w[2]), 
        .ZN(n3580) );
  INV_X1 U834 ( .A(n3581), .ZN(n8723) );
  AOI22_X1 U835 ( .A1(reg_mem[1099]), .A2(n3578), .B1(n8728), .B2(data_w[3]), 
        .ZN(n3581) );
  INV_X1 U836 ( .A(n3582), .ZN(n8724) );
  AOI22_X1 U837 ( .A1(reg_mem[1100]), .A2(n3578), .B1(n8728), .B2(data_w[4]), 
        .ZN(n3582) );
  INV_X1 U838 ( .A(n3583), .ZN(n8725) );
  AOI22_X1 U839 ( .A1(reg_mem[1101]), .A2(n3578), .B1(n8728), .B2(data_w[5]), 
        .ZN(n3583) );
  INV_X1 U840 ( .A(n3584), .ZN(n8726) );
  AOI22_X1 U841 ( .A1(reg_mem[1102]), .A2(n3578), .B1(n8728), .B2(data_w[6]), 
        .ZN(n3584) );
  INV_X1 U842 ( .A(n3585), .ZN(n8727) );
  AOI22_X1 U843 ( .A1(reg_mem[1103]), .A2(n3578), .B1(n8728), .B2(data_w[7]), 
        .ZN(n3585) );
  INV_X1 U844 ( .A(n3586), .ZN(n7567) );
  AOI22_X1 U845 ( .A1(reg_mem[1104]), .A2(n3587), .B1(n7575), .B2(data_w[0]), 
        .ZN(n3586) );
  INV_X1 U846 ( .A(n3588), .ZN(n7568) );
  AOI22_X1 U847 ( .A1(reg_mem[1105]), .A2(n3587), .B1(n7575), .B2(data_w[1]), 
        .ZN(n3588) );
  INV_X1 U848 ( .A(n3589), .ZN(n7569) );
  AOI22_X1 U849 ( .A1(reg_mem[1106]), .A2(n3587), .B1(n7575), .B2(data_w[2]), 
        .ZN(n3589) );
  INV_X1 U850 ( .A(n3590), .ZN(n7570) );
  AOI22_X1 U851 ( .A1(reg_mem[1107]), .A2(n3587), .B1(n7575), .B2(data_w[3]), 
        .ZN(n3590) );
  INV_X1 U852 ( .A(n3591), .ZN(n7571) );
  AOI22_X1 U853 ( .A1(reg_mem[1108]), .A2(n3587), .B1(n7575), .B2(data_w[4]), 
        .ZN(n3591) );
  INV_X1 U854 ( .A(n3592), .ZN(n7572) );
  AOI22_X1 U855 ( .A1(reg_mem[1109]), .A2(n3587), .B1(n7575), .B2(data_w[5]), 
        .ZN(n3592) );
  INV_X1 U856 ( .A(n3593), .ZN(n7573) );
  AOI22_X1 U857 ( .A1(reg_mem[1110]), .A2(n3587), .B1(n7575), .B2(data_w[6]), 
        .ZN(n3593) );
  INV_X1 U858 ( .A(n3594), .ZN(n7574) );
  AOI22_X1 U859 ( .A1(reg_mem[1111]), .A2(n3587), .B1(n7575), .B2(data_w[7]), 
        .ZN(n3594) );
  INV_X1 U860 ( .A(n3595), .ZN(n8144) );
  AOI22_X1 U861 ( .A1(reg_mem[1112]), .A2(n3596), .B1(n8152), .B2(data_w[0]), 
        .ZN(n3595) );
  INV_X1 U862 ( .A(n3597), .ZN(n8145) );
  AOI22_X1 U863 ( .A1(reg_mem[1113]), .A2(n3596), .B1(n8152), .B2(data_w[1]), 
        .ZN(n3597) );
  INV_X1 U864 ( .A(n3598), .ZN(n8146) );
  AOI22_X1 U865 ( .A1(reg_mem[1114]), .A2(n3596), .B1(n8152), .B2(data_w[2]), 
        .ZN(n3598) );
  INV_X1 U866 ( .A(n3599), .ZN(n8147) );
  AOI22_X1 U867 ( .A1(reg_mem[1115]), .A2(n3596), .B1(n8152), .B2(data_w[3]), 
        .ZN(n3599) );
  INV_X1 U868 ( .A(n3600), .ZN(n8148) );
  AOI22_X1 U869 ( .A1(reg_mem[1116]), .A2(n3596), .B1(n8152), .B2(data_w[4]), 
        .ZN(n3600) );
  INV_X1 U870 ( .A(n3601), .ZN(n8149) );
  AOI22_X1 U871 ( .A1(reg_mem[1117]), .A2(n3596), .B1(n8152), .B2(data_w[5]), 
        .ZN(n3601) );
  INV_X1 U872 ( .A(n3602), .ZN(n8150) );
  AOI22_X1 U873 ( .A1(reg_mem[1118]), .A2(n3596), .B1(n8152), .B2(data_w[6]), 
        .ZN(n3602) );
  INV_X1 U874 ( .A(n3603), .ZN(n8151) );
  AOI22_X1 U875 ( .A1(reg_mem[1119]), .A2(n3596), .B1(n8152), .B2(data_w[7]), 
        .ZN(n3603) );
  INV_X1 U876 ( .A(n3604), .ZN(n6847) );
  AOI22_X1 U877 ( .A1(reg_mem[1120]), .A2(n3605), .B1(n6855), .B2(data_w[0]), 
        .ZN(n3604) );
  INV_X1 U878 ( .A(n3606), .ZN(n6848) );
  AOI22_X1 U879 ( .A1(reg_mem[1121]), .A2(n3605), .B1(n6855), .B2(data_w[1]), 
        .ZN(n3606) );
  INV_X1 U880 ( .A(n3607), .ZN(n6849) );
  AOI22_X1 U881 ( .A1(reg_mem[1122]), .A2(n3605), .B1(n6855), .B2(data_w[2]), 
        .ZN(n3607) );
  INV_X1 U882 ( .A(n3608), .ZN(n6850) );
  AOI22_X1 U883 ( .A1(reg_mem[1123]), .A2(n3605), .B1(n6855), .B2(data_w[3]), 
        .ZN(n3608) );
  INV_X1 U884 ( .A(n3609), .ZN(n6851) );
  AOI22_X1 U885 ( .A1(reg_mem[1124]), .A2(n3605), .B1(n6855), .B2(data_w[4]), 
        .ZN(n3609) );
  INV_X1 U886 ( .A(n3610), .ZN(n6852) );
  AOI22_X1 U887 ( .A1(reg_mem[1125]), .A2(n3605), .B1(n6855), .B2(data_w[5]), 
        .ZN(n3610) );
  INV_X1 U888 ( .A(n3611), .ZN(n6853) );
  AOI22_X1 U889 ( .A1(reg_mem[1126]), .A2(n3605), .B1(n6855), .B2(data_w[6]), 
        .ZN(n3611) );
  INV_X1 U890 ( .A(n3612), .ZN(n6854) );
  AOI22_X1 U891 ( .A1(reg_mem[1127]), .A2(n3605), .B1(n6855), .B2(data_w[7]), 
        .ZN(n3612) );
  INV_X1 U892 ( .A(n3613), .ZN(n8576) );
  AOI22_X1 U893 ( .A1(reg_mem[1128]), .A2(n3614), .B1(n8584), .B2(data_w[0]), 
        .ZN(n3613) );
  INV_X1 U894 ( .A(n3615), .ZN(n8577) );
  AOI22_X1 U895 ( .A1(reg_mem[1129]), .A2(n3614), .B1(n8584), .B2(data_w[1]), 
        .ZN(n3615) );
  INV_X1 U896 ( .A(n3616), .ZN(n8578) );
  AOI22_X1 U897 ( .A1(reg_mem[1130]), .A2(n3614), .B1(n8584), .B2(data_w[2]), 
        .ZN(n3616) );
  INV_X1 U898 ( .A(n3617), .ZN(n8579) );
  AOI22_X1 U899 ( .A1(reg_mem[1131]), .A2(n3614), .B1(n8584), .B2(data_w[3]), 
        .ZN(n3617) );
  INV_X1 U900 ( .A(n3618), .ZN(n8580) );
  AOI22_X1 U901 ( .A1(reg_mem[1132]), .A2(n3614), .B1(n8584), .B2(data_w[4]), 
        .ZN(n3618) );
  INV_X1 U902 ( .A(n3619), .ZN(n8581) );
  AOI22_X1 U903 ( .A1(reg_mem[1133]), .A2(n3614), .B1(n8584), .B2(data_w[5]), 
        .ZN(n3619) );
  INV_X1 U904 ( .A(n3620), .ZN(n8582) );
  AOI22_X1 U905 ( .A1(reg_mem[1134]), .A2(n3614), .B1(n8584), .B2(data_w[6]), 
        .ZN(n3620) );
  INV_X1 U906 ( .A(n3621), .ZN(n8583) );
  AOI22_X1 U907 ( .A1(reg_mem[1135]), .A2(n3614), .B1(n8584), .B2(data_w[7]), 
        .ZN(n3621) );
  INV_X1 U908 ( .A(n3622), .ZN(n7423) );
  AOI22_X1 U909 ( .A1(reg_mem[1136]), .A2(n3623), .B1(n7431), .B2(data_w[0]), 
        .ZN(n3622) );
  INV_X1 U910 ( .A(n3624), .ZN(n7424) );
  AOI22_X1 U911 ( .A1(reg_mem[1137]), .A2(n3623), .B1(n7431), .B2(data_w[1]), 
        .ZN(n3624) );
  INV_X1 U912 ( .A(n3625), .ZN(n7425) );
  AOI22_X1 U913 ( .A1(reg_mem[1138]), .A2(n3623), .B1(n7431), .B2(data_w[2]), 
        .ZN(n3625) );
  INV_X1 U914 ( .A(n3626), .ZN(n7426) );
  AOI22_X1 U915 ( .A1(reg_mem[1139]), .A2(n3623), .B1(n7431), .B2(data_w[3]), 
        .ZN(n3626) );
  INV_X1 U916 ( .A(n3627), .ZN(n7427) );
  AOI22_X1 U917 ( .A1(reg_mem[1140]), .A2(n3623), .B1(n7431), .B2(data_w[4]), 
        .ZN(n3627) );
  INV_X1 U918 ( .A(n3628), .ZN(n7428) );
  AOI22_X1 U919 ( .A1(reg_mem[1141]), .A2(n3623), .B1(n7431), .B2(data_w[5]), 
        .ZN(n3628) );
  INV_X1 U920 ( .A(n3629), .ZN(n7429) );
  AOI22_X1 U921 ( .A1(reg_mem[1142]), .A2(n3623), .B1(n7431), .B2(data_w[6]), 
        .ZN(n3629) );
  INV_X1 U922 ( .A(n3630), .ZN(n7430) );
  AOI22_X1 U923 ( .A1(reg_mem[1143]), .A2(n3623), .B1(n7431), .B2(data_w[7]), 
        .ZN(n3630) );
  INV_X1 U924 ( .A(n3631), .ZN(n8000) );
  AOI22_X1 U925 ( .A1(reg_mem[1144]), .A2(n3632), .B1(n8008), .B2(data_w[0]), 
        .ZN(n3631) );
  INV_X1 U926 ( .A(n3633), .ZN(n8001) );
  AOI22_X1 U927 ( .A1(reg_mem[1145]), .A2(n3632), .B1(n8008), .B2(data_w[1]), 
        .ZN(n3633) );
  INV_X1 U928 ( .A(n3634), .ZN(n8002) );
  AOI22_X1 U929 ( .A1(reg_mem[1146]), .A2(n3632), .B1(n8008), .B2(data_w[2]), 
        .ZN(n3634) );
  INV_X1 U930 ( .A(n3635), .ZN(n8003) );
  AOI22_X1 U931 ( .A1(reg_mem[1147]), .A2(n3632), .B1(n8008), .B2(data_w[3]), 
        .ZN(n3635) );
  INV_X1 U932 ( .A(n3636), .ZN(n8004) );
  AOI22_X1 U933 ( .A1(reg_mem[1148]), .A2(n3632), .B1(n8008), .B2(data_w[4]), 
        .ZN(n3636) );
  INV_X1 U934 ( .A(n3637), .ZN(n8005) );
  AOI22_X1 U935 ( .A1(reg_mem[1149]), .A2(n3632), .B1(n8008), .B2(data_w[5]), 
        .ZN(n3637) );
  INV_X1 U936 ( .A(n3638), .ZN(n8006) );
  AOI22_X1 U937 ( .A1(reg_mem[1150]), .A2(n3632), .B1(n8008), .B2(data_w[6]), 
        .ZN(n3638) );
  INV_X1 U938 ( .A(n3639), .ZN(n8007) );
  AOI22_X1 U939 ( .A1(reg_mem[1151]), .A2(n3632), .B1(n8008), .B2(data_w[7]), 
        .ZN(n3639) );
  INV_X1 U940 ( .A(n3641), .ZN(n7270) );
  AOI22_X1 U941 ( .A1(reg_mem[1152]), .A2(n3642), .B1(n7278), .B2(data_w[0]), 
        .ZN(n3641) );
  INV_X1 U942 ( .A(n3643), .ZN(n7271) );
  AOI22_X1 U943 ( .A1(reg_mem[1153]), .A2(n3642), .B1(n7278), .B2(data_w[1]), 
        .ZN(n3643) );
  INV_X1 U944 ( .A(n3644), .ZN(n7272) );
  AOI22_X1 U945 ( .A1(reg_mem[1154]), .A2(n3642), .B1(n7278), .B2(data_w[2]), 
        .ZN(n3644) );
  INV_X1 U946 ( .A(n3645), .ZN(n7273) );
  AOI22_X1 U947 ( .A1(reg_mem[1155]), .A2(n3642), .B1(n7278), .B2(data_w[3]), 
        .ZN(n3645) );
  INV_X1 U948 ( .A(n3646), .ZN(n7274) );
  AOI22_X1 U949 ( .A1(reg_mem[1156]), .A2(n3642), .B1(n7278), .B2(data_w[4]), 
        .ZN(n3646) );
  INV_X1 U950 ( .A(n3647), .ZN(n7275) );
  AOI22_X1 U951 ( .A1(reg_mem[1157]), .A2(n3642), .B1(n7278), .B2(data_w[5]), 
        .ZN(n3647) );
  INV_X1 U952 ( .A(n3648), .ZN(n7276) );
  AOI22_X1 U953 ( .A1(reg_mem[1158]), .A2(n3642), .B1(n7278), .B2(data_w[6]), 
        .ZN(n3648) );
  INV_X1 U954 ( .A(n3649), .ZN(n7277) );
  AOI22_X1 U955 ( .A1(reg_mem[1159]), .A2(n3642), .B1(n7278), .B2(data_w[7]), 
        .ZN(n3649) );
  INV_X1 U956 ( .A(n3651), .ZN(n8999) );
  AOI22_X1 U957 ( .A1(reg_mem[1160]), .A2(n3652), .B1(n9007), .B2(data_w[0]), 
        .ZN(n3651) );
  INV_X1 U958 ( .A(n3653), .ZN(n9000) );
  AOI22_X1 U959 ( .A1(reg_mem[1161]), .A2(n3652), .B1(n9007), .B2(data_w[1]), 
        .ZN(n3653) );
  INV_X1 U960 ( .A(n3654), .ZN(n9001) );
  AOI22_X1 U961 ( .A1(reg_mem[1162]), .A2(n3652), .B1(n9007), .B2(data_w[2]), 
        .ZN(n3654) );
  INV_X1 U962 ( .A(n3655), .ZN(n9002) );
  AOI22_X1 U963 ( .A1(reg_mem[1163]), .A2(n3652), .B1(n9007), .B2(data_w[3]), 
        .ZN(n3655) );
  INV_X1 U964 ( .A(n3656), .ZN(n9003) );
  AOI22_X1 U965 ( .A1(reg_mem[1164]), .A2(n3652), .B1(n9007), .B2(data_w[4]), 
        .ZN(n3656) );
  INV_X1 U966 ( .A(n3657), .ZN(n9004) );
  AOI22_X1 U967 ( .A1(reg_mem[1165]), .A2(n3652), .B1(n9007), .B2(data_w[5]), 
        .ZN(n3657) );
  INV_X1 U968 ( .A(n3658), .ZN(n9005) );
  AOI22_X1 U969 ( .A1(reg_mem[1166]), .A2(n3652), .B1(n9007), .B2(data_w[6]), 
        .ZN(n3658) );
  INV_X1 U970 ( .A(n3659), .ZN(n9006) );
  AOI22_X1 U971 ( .A1(reg_mem[1167]), .A2(n3652), .B1(n9007), .B2(data_w[7]), 
        .ZN(n3659) );
  INV_X1 U972 ( .A(n3660), .ZN(n7846) );
  AOI22_X1 U973 ( .A1(reg_mem[1168]), .A2(n3661), .B1(n7854), .B2(data_w[0]), 
        .ZN(n3660) );
  INV_X1 U974 ( .A(n3662), .ZN(n7847) );
  AOI22_X1 U975 ( .A1(reg_mem[1169]), .A2(n3661), .B1(n7854), .B2(data_w[1]), 
        .ZN(n3662) );
  INV_X1 U976 ( .A(n3663), .ZN(n7848) );
  AOI22_X1 U977 ( .A1(reg_mem[1170]), .A2(n3661), .B1(n7854), .B2(data_w[2]), 
        .ZN(n3663) );
  INV_X1 U978 ( .A(n3664), .ZN(n7849) );
  AOI22_X1 U979 ( .A1(reg_mem[1171]), .A2(n3661), .B1(n7854), .B2(data_w[3]), 
        .ZN(n3664) );
  INV_X1 U980 ( .A(n3665), .ZN(n7850) );
  AOI22_X1 U981 ( .A1(reg_mem[1172]), .A2(n3661), .B1(n7854), .B2(data_w[4]), 
        .ZN(n3665) );
  INV_X1 U982 ( .A(n3666), .ZN(n7851) );
  AOI22_X1 U983 ( .A1(reg_mem[1173]), .A2(n3661), .B1(n7854), .B2(data_w[5]), 
        .ZN(n3666) );
  INV_X1 U984 ( .A(n3667), .ZN(n7852) );
  AOI22_X1 U985 ( .A1(reg_mem[1174]), .A2(n3661), .B1(n7854), .B2(data_w[6]), 
        .ZN(n3667) );
  INV_X1 U986 ( .A(n3668), .ZN(n7853) );
  AOI22_X1 U987 ( .A1(reg_mem[1175]), .A2(n3661), .B1(n7854), .B2(data_w[7]), 
        .ZN(n3668) );
  INV_X1 U988 ( .A(n3669), .ZN(n8423) );
  AOI22_X1 U989 ( .A1(reg_mem[1176]), .A2(n3670), .B1(n8431), .B2(data_w[0]), 
        .ZN(n3669) );
  INV_X1 U990 ( .A(n3671), .ZN(n8424) );
  AOI22_X1 U991 ( .A1(reg_mem[1177]), .A2(n3670), .B1(n8431), .B2(data_w[1]), 
        .ZN(n3671) );
  INV_X1 U992 ( .A(n3672), .ZN(n8425) );
  AOI22_X1 U993 ( .A1(reg_mem[1178]), .A2(n3670), .B1(n8431), .B2(data_w[2]), 
        .ZN(n3672) );
  INV_X1 U994 ( .A(n3673), .ZN(n8426) );
  AOI22_X1 U995 ( .A1(reg_mem[1179]), .A2(n3670), .B1(n8431), .B2(data_w[3]), 
        .ZN(n3673) );
  INV_X1 U996 ( .A(n3674), .ZN(n8427) );
  AOI22_X1 U997 ( .A1(reg_mem[1180]), .A2(n3670), .B1(n8431), .B2(data_w[4]), 
        .ZN(n3674) );
  INV_X1 U998 ( .A(n3675), .ZN(n8428) );
  AOI22_X1 U999 ( .A1(reg_mem[1181]), .A2(n3670), .B1(n8431), .B2(data_w[5]), 
        .ZN(n3675) );
  INV_X1 U1000 ( .A(n3676), .ZN(n8429) );
  AOI22_X1 U1001 ( .A1(reg_mem[1182]), .A2(n3670), .B1(n8431), .B2(data_w[6]), 
        .ZN(n3676) );
  INV_X1 U1002 ( .A(n3677), .ZN(n8430) );
  AOI22_X1 U1003 ( .A1(reg_mem[1183]), .A2(n3670), .B1(n8431), .B2(data_w[7]), 
        .ZN(n3677) );
  INV_X1 U1004 ( .A(n3678), .ZN(n7126) );
  AOI22_X1 U1005 ( .A1(reg_mem[1184]), .A2(n3679), .B1(n7134), .B2(data_w[0]), 
        .ZN(n3678) );
  INV_X1 U1006 ( .A(n3680), .ZN(n7127) );
  AOI22_X1 U1007 ( .A1(reg_mem[1185]), .A2(n3679), .B1(n7134), .B2(data_w[1]), 
        .ZN(n3680) );
  INV_X1 U1008 ( .A(n3681), .ZN(n7128) );
  AOI22_X1 U1009 ( .A1(reg_mem[1186]), .A2(n3679), .B1(n7134), .B2(data_w[2]), 
        .ZN(n3681) );
  INV_X1 U1010 ( .A(n3682), .ZN(n7129) );
  AOI22_X1 U1011 ( .A1(reg_mem[1187]), .A2(n3679), .B1(n7134), .B2(data_w[3]), 
        .ZN(n3682) );
  INV_X1 U1012 ( .A(n3683), .ZN(n7130) );
  AOI22_X1 U1013 ( .A1(reg_mem[1188]), .A2(n3679), .B1(n7134), .B2(data_w[4]), 
        .ZN(n3683) );
  INV_X1 U1014 ( .A(n3684), .ZN(n7131) );
  AOI22_X1 U1015 ( .A1(reg_mem[1189]), .A2(n3679), .B1(n7134), .B2(data_w[5]), 
        .ZN(n3684) );
  INV_X1 U1016 ( .A(n3685), .ZN(n7132) );
  AOI22_X1 U1017 ( .A1(reg_mem[1190]), .A2(n3679), .B1(n7134), .B2(data_w[6]), 
        .ZN(n3685) );
  INV_X1 U1018 ( .A(n3686), .ZN(n7133) );
  AOI22_X1 U1019 ( .A1(reg_mem[1191]), .A2(n3679), .B1(n7134), .B2(data_w[7]), 
        .ZN(n3686) );
  INV_X1 U1020 ( .A(n3687), .ZN(n8855) );
  AOI22_X1 U1021 ( .A1(reg_mem[1192]), .A2(n3688), .B1(n8863), .B2(data_w[0]), 
        .ZN(n3687) );
  INV_X1 U1022 ( .A(n3689), .ZN(n8856) );
  AOI22_X1 U1023 ( .A1(reg_mem[1193]), .A2(n3688), .B1(n8863), .B2(data_w[1]), 
        .ZN(n3689) );
  INV_X1 U1024 ( .A(n3690), .ZN(n8857) );
  AOI22_X1 U1025 ( .A1(reg_mem[1194]), .A2(n3688), .B1(n8863), .B2(data_w[2]), 
        .ZN(n3690) );
  INV_X1 U1026 ( .A(n3691), .ZN(n8858) );
  AOI22_X1 U1027 ( .A1(reg_mem[1195]), .A2(n3688), .B1(n8863), .B2(data_w[3]), 
        .ZN(n3691) );
  INV_X1 U1028 ( .A(n3692), .ZN(n8859) );
  AOI22_X1 U1029 ( .A1(reg_mem[1196]), .A2(n3688), .B1(n8863), .B2(data_w[4]), 
        .ZN(n3692) );
  INV_X1 U1030 ( .A(n3693), .ZN(n8860) );
  AOI22_X1 U1031 ( .A1(reg_mem[1197]), .A2(n3688), .B1(n8863), .B2(data_w[5]), 
        .ZN(n3693) );
  INV_X1 U1032 ( .A(n3694), .ZN(n8861) );
  AOI22_X1 U1033 ( .A1(reg_mem[1198]), .A2(n3688), .B1(n8863), .B2(data_w[6]), 
        .ZN(n3694) );
  INV_X1 U1034 ( .A(n3695), .ZN(n8862) );
  AOI22_X1 U1035 ( .A1(reg_mem[1199]), .A2(n3688), .B1(n8863), .B2(data_w[7]), 
        .ZN(n3695) );
  INV_X1 U1036 ( .A(n3696), .ZN(n7702) );
  AOI22_X1 U1037 ( .A1(reg_mem[1200]), .A2(n3697), .B1(n7710), .B2(data_w[0]), 
        .ZN(n3696) );
  INV_X1 U1038 ( .A(n3698), .ZN(n7703) );
  AOI22_X1 U1039 ( .A1(reg_mem[1201]), .A2(n3697), .B1(n7710), .B2(data_w[1]), 
        .ZN(n3698) );
  INV_X1 U1040 ( .A(n3699), .ZN(n7704) );
  AOI22_X1 U1041 ( .A1(reg_mem[1202]), .A2(n3697), .B1(n7710), .B2(data_w[2]), 
        .ZN(n3699) );
  INV_X1 U1042 ( .A(n3700), .ZN(n7705) );
  AOI22_X1 U1043 ( .A1(reg_mem[1203]), .A2(n3697), .B1(n7710), .B2(data_w[3]), 
        .ZN(n3700) );
  INV_X1 U1044 ( .A(n3701), .ZN(n7706) );
  AOI22_X1 U1045 ( .A1(reg_mem[1204]), .A2(n3697), .B1(n7710), .B2(data_w[4]), 
        .ZN(n3701) );
  INV_X1 U1046 ( .A(n3702), .ZN(n7707) );
  AOI22_X1 U1047 ( .A1(reg_mem[1205]), .A2(n3697), .B1(n7710), .B2(data_w[5]), 
        .ZN(n3702) );
  INV_X1 U1048 ( .A(n3703), .ZN(n7708) );
  AOI22_X1 U1049 ( .A1(reg_mem[1206]), .A2(n3697), .B1(n7710), .B2(data_w[6]), 
        .ZN(n3703) );
  INV_X1 U1050 ( .A(n3704), .ZN(n7709) );
  AOI22_X1 U1051 ( .A1(reg_mem[1207]), .A2(n3697), .B1(n7710), .B2(data_w[7]), 
        .ZN(n3704) );
  INV_X1 U1052 ( .A(n3705), .ZN(n8279) );
  AOI22_X1 U1053 ( .A1(reg_mem[1208]), .A2(n3706), .B1(n8287), .B2(data_w[0]), 
        .ZN(n3705) );
  INV_X1 U1054 ( .A(n3707), .ZN(n8280) );
  AOI22_X1 U1055 ( .A1(reg_mem[1209]), .A2(n3706), .B1(n8287), .B2(data_w[1]), 
        .ZN(n3707) );
  INV_X1 U1056 ( .A(n3708), .ZN(n8281) );
  AOI22_X1 U1057 ( .A1(reg_mem[1210]), .A2(n3706), .B1(n8287), .B2(data_w[2]), 
        .ZN(n3708) );
  INV_X1 U1058 ( .A(n3709), .ZN(n8282) );
  AOI22_X1 U1059 ( .A1(reg_mem[1211]), .A2(n3706), .B1(n8287), .B2(data_w[3]), 
        .ZN(n3709) );
  INV_X1 U1060 ( .A(n3710), .ZN(n8283) );
  AOI22_X1 U1061 ( .A1(reg_mem[1212]), .A2(n3706), .B1(n8287), .B2(data_w[4]), 
        .ZN(n3710) );
  INV_X1 U1062 ( .A(n3711), .ZN(n8284) );
  AOI22_X1 U1063 ( .A1(reg_mem[1213]), .A2(n3706), .B1(n8287), .B2(data_w[5]), 
        .ZN(n3711) );
  INV_X1 U1064 ( .A(n3712), .ZN(n8285) );
  AOI22_X1 U1065 ( .A1(reg_mem[1214]), .A2(n3706), .B1(n8287), .B2(data_w[6]), 
        .ZN(n3712) );
  INV_X1 U1066 ( .A(n3713), .ZN(n8286) );
  AOI22_X1 U1067 ( .A1(reg_mem[1215]), .A2(n3706), .B1(n8287), .B2(data_w[7]), 
        .ZN(n3713) );
  INV_X1 U1068 ( .A(n3714), .ZN(n6982) );
  AOI22_X1 U1069 ( .A1(reg_mem[1216]), .A2(n3715), .B1(n6990), .B2(data_w[0]), 
        .ZN(n3714) );
  INV_X1 U1070 ( .A(n3716), .ZN(n6983) );
  AOI22_X1 U1071 ( .A1(reg_mem[1217]), .A2(n3715), .B1(n6990), .B2(data_w[1]), 
        .ZN(n3716) );
  INV_X1 U1072 ( .A(n3717), .ZN(n6984) );
  AOI22_X1 U1073 ( .A1(reg_mem[1218]), .A2(n3715), .B1(n6990), .B2(data_w[2]), 
        .ZN(n3717) );
  INV_X1 U1074 ( .A(n3718), .ZN(n6985) );
  AOI22_X1 U1075 ( .A1(reg_mem[1219]), .A2(n3715), .B1(n6990), .B2(data_w[3]), 
        .ZN(n3718) );
  INV_X1 U1076 ( .A(n3719), .ZN(n6986) );
  AOI22_X1 U1077 ( .A1(reg_mem[1220]), .A2(n3715), .B1(n6990), .B2(data_w[4]), 
        .ZN(n3719) );
  INV_X1 U1078 ( .A(n3720), .ZN(n6987) );
  AOI22_X1 U1079 ( .A1(reg_mem[1221]), .A2(n3715), .B1(n6990), .B2(data_w[5]), 
        .ZN(n3720) );
  INV_X1 U1080 ( .A(n3721), .ZN(n6988) );
  AOI22_X1 U1081 ( .A1(reg_mem[1222]), .A2(n3715), .B1(n6990), .B2(data_w[6]), 
        .ZN(n3721) );
  INV_X1 U1082 ( .A(n3722), .ZN(n6989) );
  AOI22_X1 U1083 ( .A1(reg_mem[1223]), .A2(n3715), .B1(n6990), .B2(data_w[7]), 
        .ZN(n3722) );
  INV_X1 U1084 ( .A(n3723), .ZN(n8711) );
  AOI22_X1 U1085 ( .A1(reg_mem[1224]), .A2(n3724), .B1(n8719), .B2(data_w[0]), 
        .ZN(n3723) );
  INV_X1 U1086 ( .A(n3725), .ZN(n8712) );
  AOI22_X1 U1087 ( .A1(reg_mem[1225]), .A2(n3724), .B1(n8719), .B2(data_w[1]), 
        .ZN(n3725) );
  INV_X1 U1088 ( .A(n3726), .ZN(n8713) );
  AOI22_X1 U1089 ( .A1(reg_mem[1226]), .A2(n3724), .B1(n8719), .B2(data_w[2]), 
        .ZN(n3726) );
  INV_X1 U1090 ( .A(n3727), .ZN(n8714) );
  AOI22_X1 U1091 ( .A1(reg_mem[1227]), .A2(n3724), .B1(n8719), .B2(data_w[3]), 
        .ZN(n3727) );
  INV_X1 U1092 ( .A(n3728), .ZN(n8715) );
  AOI22_X1 U1093 ( .A1(reg_mem[1228]), .A2(n3724), .B1(n8719), .B2(data_w[4]), 
        .ZN(n3728) );
  INV_X1 U1094 ( .A(n3729), .ZN(n8716) );
  AOI22_X1 U1095 ( .A1(reg_mem[1229]), .A2(n3724), .B1(n8719), .B2(data_w[5]), 
        .ZN(n3729) );
  INV_X1 U1096 ( .A(n3730), .ZN(n8717) );
  AOI22_X1 U1097 ( .A1(reg_mem[1230]), .A2(n3724), .B1(n8719), .B2(data_w[6]), 
        .ZN(n3730) );
  INV_X1 U1098 ( .A(n3731), .ZN(n8718) );
  AOI22_X1 U1099 ( .A1(reg_mem[1231]), .A2(n3724), .B1(n8719), .B2(data_w[7]), 
        .ZN(n3731) );
  INV_X1 U1100 ( .A(n3732), .ZN(n7558) );
  AOI22_X1 U1101 ( .A1(reg_mem[1232]), .A2(n3733), .B1(n7566), .B2(data_w[0]), 
        .ZN(n3732) );
  INV_X1 U1102 ( .A(n3734), .ZN(n7559) );
  AOI22_X1 U1103 ( .A1(reg_mem[1233]), .A2(n3733), .B1(n7566), .B2(data_w[1]), 
        .ZN(n3734) );
  INV_X1 U1104 ( .A(n3735), .ZN(n7560) );
  AOI22_X1 U1105 ( .A1(reg_mem[1234]), .A2(n3733), .B1(n7566), .B2(data_w[2]), 
        .ZN(n3735) );
  INV_X1 U1106 ( .A(n3736), .ZN(n7561) );
  AOI22_X1 U1107 ( .A1(reg_mem[1235]), .A2(n3733), .B1(n7566), .B2(data_w[3]), 
        .ZN(n3736) );
  INV_X1 U1108 ( .A(n3737), .ZN(n7562) );
  AOI22_X1 U1109 ( .A1(reg_mem[1236]), .A2(n3733), .B1(n7566), .B2(data_w[4]), 
        .ZN(n3737) );
  INV_X1 U1110 ( .A(n3738), .ZN(n7563) );
  AOI22_X1 U1111 ( .A1(reg_mem[1237]), .A2(n3733), .B1(n7566), .B2(data_w[5]), 
        .ZN(n3738) );
  INV_X1 U1112 ( .A(n3739), .ZN(n7564) );
  AOI22_X1 U1113 ( .A1(reg_mem[1238]), .A2(n3733), .B1(n7566), .B2(data_w[6]), 
        .ZN(n3739) );
  INV_X1 U1114 ( .A(n3740), .ZN(n7565) );
  AOI22_X1 U1115 ( .A1(reg_mem[1239]), .A2(n3733), .B1(n7566), .B2(data_w[7]), 
        .ZN(n3740) );
  INV_X1 U1116 ( .A(n3741), .ZN(n8135) );
  AOI22_X1 U1117 ( .A1(reg_mem[1240]), .A2(n3742), .B1(n8143), .B2(data_w[0]), 
        .ZN(n3741) );
  INV_X1 U1118 ( .A(n3743), .ZN(n8136) );
  AOI22_X1 U1119 ( .A1(reg_mem[1241]), .A2(n3742), .B1(n8143), .B2(data_w[1]), 
        .ZN(n3743) );
  INV_X1 U1120 ( .A(n3744), .ZN(n8137) );
  AOI22_X1 U1121 ( .A1(reg_mem[1242]), .A2(n3742), .B1(n8143), .B2(data_w[2]), 
        .ZN(n3744) );
  INV_X1 U1122 ( .A(n3745), .ZN(n8138) );
  AOI22_X1 U1123 ( .A1(reg_mem[1243]), .A2(n3742), .B1(n8143), .B2(data_w[3]), 
        .ZN(n3745) );
  INV_X1 U1124 ( .A(n3746), .ZN(n8139) );
  AOI22_X1 U1125 ( .A1(reg_mem[1244]), .A2(n3742), .B1(n8143), .B2(data_w[4]), 
        .ZN(n3746) );
  INV_X1 U1126 ( .A(n3747), .ZN(n8140) );
  AOI22_X1 U1127 ( .A1(reg_mem[1245]), .A2(n3742), .B1(n8143), .B2(data_w[5]), 
        .ZN(n3747) );
  INV_X1 U1128 ( .A(n3748), .ZN(n8141) );
  AOI22_X1 U1129 ( .A1(reg_mem[1246]), .A2(n3742), .B1(n8143), .B2(data_w[6]), 
        .ZN(n3748) );
  INV_X1 U1130 ( .A(n3749), .ZN(n8142) );
  AOI22_X1 U1131 ( .A1(reg_mem[1247]), .A2(n3742), .B1(n8143), .B2(data_w[7]), 
        .ZN(n3749) );
  INV_X1 U1132 ( .A(n3750), .ZN(n6838) );
  AOI22_X1 U1133 ( .A1(reg_mem[1248]), .A2(n3751), .B1(n6846), .B2(data_w[0]), 
        .ZN(n3750) );
  INV_X1 U1134 ( .A(n3752), .ZN(n6839) );
  AOI22_X1 U1135 ( .A1(reg_mem[1249]), .A2(n3751), .B1(n6846), .B2(data_w[1]), 
        .ZN(n3752) );
  INV_X1 U1136 ( .A(n3753), .ZN(n6840) );
  AOI22_X1 U1137 ( .A1(reg_mem[1250]), .A2(n3751), .B1(n6846), .B2(data_w[2]), 
        .ZN(n3753) );
  INV_X1 U1138 ( .A(n3754), .ZN(n6841) );
  AOI22_X1 U1139 ( .A1(reg_mem[1251]), .A2(n3751), .B1(n6846), .B2(data_w[3]), 
        .ZN(n3754) );
  INV_X1 U1140 ( .A(n3755), .ZN(n6842) );
  AOI22_X1 U1141 ( .A1(reg_mem[1252]), .A2(n3751), .B1(n6846), .B2(data_w[4]), 
        .ZN(n3755) );
  INV_X1 U1142 ( .A(n3756), .ZN(n6843) );
  AOI22_X1 U1143 ( .A1(reg_mem[1253]), .A2(n3751), .B1(n6846), .B2(data_w[5]), 
        .ZN(n3756) );
  INV_X1 U1144 ( .A(n3757), .ZN(n6844) );
  AOI22_X1 U1145 ( .A1(reg_mem[1254]), .A2(n3751), .B1(n6846), .B2(data_w[6]), 
        .ZN(n3757) );
  INV_X1 U1146 ( .A(n3758), .ZN(n6845) );
  AOI22_X1 U1147 ( .A1(reg_mem[1255]), .A2(n3751), .B1(n6846), .B2(data_w[7]), 
        .ZN(n3758) );
  INV_X1 U1148 ( .A(n3759), .ZN(n8567) );
  AOI22_X1 U1149 ( .A1(reg_mem[1256]), .A2(n3760), .B1(n8575), .B2(data_w[0]), 
        .ZN(n3759) );
  INV_X1 U1150 ( .A(n3761), .ZN(n8568) );
  AOI22_X1 U1151 ( .A1(reg_mem[1257]), .A2(n3760), .B1(n8575), .B2(data_w[1]), 
        .ZN(n3761) );
  INV_X1 U1152 ( .A(n3762), .ZN(n8569) );
  AOI22_X1 U1153 ( .A1(reg_mem[1258]), .A2(n3760), .B1(n8575), .B2(data_w[2]), 
        .ZN(n3762) );
  INV_X1 U1154 ( .A(n3763), .ZN(n8570) );
  AOI22_X1 U1155 ( .A1(reg_mem[1259]), .A2(n3760), .B1(n8575), .B2(data_w[3]), 
        .ZN(n3763) );
  INV_X1 U1156 ( .A(n3764), .ZN(n8571) );
  AOI22_X1 U1157 ( .A1(reg_mem[1260]), .A2(n3760), .B1(n8575), .B2(data_w[4]), 
        .ZN(n3764) );
  INV_X1 U1158 ( .A(n3765), .ZN(n8572) );
  AOI22_X1 U1159 ( .A1(reg_mem[1261]), .A2(n3760), .B1(n8575), .B2(data_w[5]), 
        .ZN(n3765) );
  INV_X1 U1160 ( .A(n3766), .ZN(n8573) );
  AOI22_X1 U1161 ( .A1(reg_mem[1262]), .A2(n3760), .B1(n8575), .B2(data_w[6]), 
        .ZN(n3766) );
  INV_X1 U1162 ( .A(n3767), .ZN(n8574) );
  AOI22_X1 U1163 ( .A1(reg_mem[1263]), .A2(n3760), .B1(n8575), .B2(data_w[7]), 
        .ZN(n3767) );
  INV_X1 U1164 ( .A(n3768), .ZN(n7414) );
  AOI22_X1 U1165 ( .A1(reg_mem[1264]), .A2(n3769), .B1(n7422), .B2(data_w[0]), 
        .ZN(n3768) );
  INV_X1 U1166 ( .A(n3770), .ZN(n7415) );
  AOI22_X1 U1167 ( .A1(reg_mem[1265]), .A2(n3769), .B1(n7422), .B2(data_w[1]), 
        .ZN(n3770) );
  INV_X1 U1168 ( .A(n3771), .ZN(n7416) );
  AOI22_X1 U1169 ( .A1(reg_mem[1266]), .A2(n3769), .B1(n7422), .B2(data_w[2]), 
        .ZN(n3771) );
  INV_X1 U1170 ( .A(n3772), .ZN(n7417) );
  AOI22_X1 U1171 ( .A1(reg_mem[1267]), .A2(n3769), .B1(n7422), .B2(data_w[3]), 
        .ZN(n3772) );
  INV_X1 U1172 ( .A(n3773), .ZN(n7418) );
  AOI22_X1 U1173 ( .A1(reg_mem[1268]), .A2(n3769), .B1(n7422), .B2(data_w[4]), 
        .ZN(n3773) );
  INV_X1 U1174 ( .A(n3774), .ZN(n7419) );
  AOI22_X1 U1175 ( .A1(reg_mem[1269]), .A2(n3769), .B1(n7422), .B2(data_w[5]), 
        .ZN(n3774) );
  INV_X1 U1176 ( .A(n3775), .ZN(n7420) );
  AOI22_X1 U1177 ( .A1(reg_mem[1270]), .A2(n3769), .B1(n7422), .B2(data_w[6]), 
        .ZN(n3775) );
  INV_X1 U1178 ( .A(n3776), .ZN(n7421) );
  AOI22_X1 U1179 ( .A1(reg_mem[1271]), .A2(n3769), .B1(n7422), .B2(data_w[7]), 
        .ZN(n3776) );
  INV_X1 U1180 ( .A(n3777), .ZN(n7991) );
  AOI22_X1 U1181 ( .A1(reg_mem[1272]), .A2(n3778), .B1(n7999), .B2(data_w[0]), 
        .ZN(n3777) );
  INV_X1 U1182 ( .A(n3779), .ZN(n7992) );
  AOI22_X1 U1183 ( .A1(reg_mem[1273]), .A2(n3778), .B1(n7999), .B2(data_w[1]), 
        .ZN(n3779) );
  INV_X1 U1184 ( .A(n3780), .ZN(n7993) );
  AOI22_X1 U1185 ( .A1(reg_mem[1274]), .A2(n3778), .B1(n7999), .B2(data_w[2]), 
        .ZN(n3780) );
  INV_X1 U1186 ( .A(n3781), .ZN(n7994) );
  AOI22_X1 U1187 ( .A1(reg_mem[1275]), .A2(n3778), .B1(n7999), .B2(data_w[3]), 
        .ZN(n3781) );
  INV_X1 U1188 ( .A(n3782), .ZN(n7995) );
  AOI22_X1 U1189 ( .A1(reg_mem[1276]), .A2(n3778), .B1(n7999), .B2(data_w[4]), 
        .ZN(n3782) );
  INV_X1 U1190 ( .A(n3783), .ZN(n7996) );
  AOI22_X1 U1191 ( .A1(reg_mem[1277]), .A2(n3778), .B1(n7999), .B2(data_w[5]), 
        .ZN(n3783) );
  INV_X1 U1192 ( .A(n3784), .ZN(n7997) );
  AOI22_X1 U1193 ( .A1(reg_mem[1278]), .A2(n3778), .B1(n7999), .B2(data_w[6]), 
        .ZN(n3784) );
  INV_X1 U1194 ( .A(n3785), .ZN(n7998) );
  AOI22_X1 U1195 ( .A1(reg_mem[1279]), .A2(n3778), .B1(n7999), .B2(data_w[7]), 
        .ZN(n3785) );
  INV_X1 U1196 ( .A(n3786), .ZN(n7261) );
  AOI22_X1 U1197 ( .A1(reg_mem[1280]), .A2(n3787), .B1(n7269), .B2(data_w[0]), 
        .ZN(n3786) );
  INV_X1 U1198 ( .A(n3788), .ZN(n7262) );
  AOI22_X1 U1199 ( .A1(reg_mem[1281]), .A2(n3787), .B1(n7269), .B2(data_w[1]), 
        .ZN(n3788) );
  INV_X1 U1200 ( .A(n3789), .ZN(n7263) );
  AOI22_X1 U1201 ( .A1(reg_mem[1282]), .A2(n3787), .B1(n7269), .B2(data_w[2]), 
        .ZN(n3789) );
  INV_X1 U1202 ( .A(n3790), .ZN(n7264) );
  AOI22_X1 U1203 ( .A1(reg_mem[1283]), .A2(n3787), .B1(n7269), .B2(data_w[3]), 
        .ZN(n3790) );
  INV_X1 U1204 ( .A(n3791), .ZN(n7265) );
  AOI22_X1 U1205 ( .A1(reg_mem[1284]), .A2(n3787), .B1(n7269), .B2(data_w[4]), 
        .ZN(n3791) );
  INV_X1 U1206 ( .A(n3792), .ZN(n7266) );
  AOI22_X1 U1207 ( .A1(reg_mem[1285]), .A2(n3787), .B1(n7269), .B2(data_w[5]), 
        .ZN(n3792) );
  INV_X1 U1208 ( .A(n3793), .ZN(n7267) );
  AOI22_X1 U1209 ( .A1(reg_mem[1286]), .A2(n3787), .B1(n7269), .B2(data_w[6]), 
        .ZN(n3793) );
  INV_X1 U1210 ( .A(n3794), .ZN(n7268) );
  AOI22_X1 U1211 ( .A1(reg_mem[1287]), .A2(n3787), .B1(n7269), .B2(data_w[7]), 
        .ZN(n3794) );
  INV_X1 U1212 ( .A(n3796), .ZN(n8990) );
  AOI22_X1 U1213 ( .A1(reg_mem[1288]), .A2(n3797), .B1(n8998), .B2(data_w[0]), 
        .ZN(n3796) );
  INV_X1 U1214 ( .A(n3798), .ZN(n8991) );
  AOI22_X1 U1215 ( .A1(reg_mem[1289]), .A2(n3797), .B1(n8998), .B2(data_w[1]), 
        .ZN(n3798) );
  INV_X1 U1216 ( .A(n3799), .ZN(n8992) );
  AOI22_X1 U1217 ( .A1(reg_mem[1290]), .A2(n3797), .B1(n8998), .B2(data_w[2]), 
        .ZN(n3799) );
  INV_X1 U1218 ( .A(n3800), .ZN(n8993) );
  AOI22_X1 U1219 ( .A1(reg_mem[1291]), .A2(n3797), .B1(n8998), .B2(data_w[3]), 
        .ZN(n3800) );
  INV_X1 U1220 ( .A(n3801), .ZN(n8994) );
  AOI22_X1 U1221 ( .A1(reg_mem[1292]), .A2(n3797), .B1(n8998), .B2(data_w[4]), 
        .ZN(n3801) );
  INV_X1 U1222 ( .A(n3802), .ZN(n8995) );
  AOI22_X1 U1223 ( .A1(reg_mem[1293]), .A2(n3797), .B1(n8998), .B2(data_w[5]), 
        .ZN(n3802) );
  INV_X1 U1224 ( .A(n3803), .ZN(n8996) );
  AOI22_X1 U1225 ( .A1(reg_mem[1294]), .A2(n3797), .B1(n8998), .B2(data_w[6]), 
        .ZN(n3803) );
  INV_X1 U1226 ( .A(n3804), .ZN(n8997) );
  AOI22_X1 U1227 ( .A1(reg_mem[1295]), .A2(n3797), .B1(n8998), .B2(data_w[7]), 
        .ZN(n3804) );
  INV_X1 U1228 ( .A(n3805), .ZN(n7837) );
  AOI22_X1 U1229 ( .A1(reg_mem[1296]), .A2(n3806), .B1(n7845), .B2(data_w[0]), 
        .ZN(n3805) );
  INV_X1 U1230 ( .A(n3807), .ZN(n7838) );
  AOI22_X1 U1231 ( .A1(reg_mem[1297]), .A2(n3806), .B1(n7845), .B2(data_w[1]), 
        .ZN(n3807) );
  INV_X1 U1232 ( .A(n3808), .ZN(n7839) );
  AOI22_X1 U1233 ( .A1(reg_mem[1298]), .A2(n3806), .B1(n7845), .B2(data_w[2]), 
        .ZN(n3808) );
  INV_X1 U1234 ( .A(n3809), .ZN(n7840) );
  AOI22_X1 U1235 ( .A1(reg_mem[1299]), .A2(n3806), .B1(n7845), .B2(data_w[3]), 
        .ZN(n3809) );
  INV_X1 U1236 ( .A(n3810), .ZN(n7841) );
  AOI22_X1 U1237 ( .A1(reg_mem[1300]), .A2(n3806), .B1(n7845), .B2(data_w[4]), 
        .ZN(n3810) );
  INV_X1 U1238 ( .A(n3811), .ZN(n7842) );
  AOI22_X1 U1239 ( .A1(reg_mem[1301]), .A2(n3806), .B1(n7845), .B2(data_w[5]), 
        .ZN(n3811) );
  INV_X1 U1240 ( .A(n3812), .ZN(n7843) );
  AOI22_X1 U1241 ( .A1(reg_mem[1302]), .A2(n3806), .B1(n7845), .B2(data_w[6]), 
        .ZN(n3812) );
  INV_X1 U1242 ( .A(n3813), .ZN(n7844) );
  AOI22_X1 U1243 ( .A1(reg_mem[1303]), .A2(n3806), .B1(n7845), .B2(data_w[7]), 
        .ZN(n3813) );
  INV_X1 U1244 ( .A(n3814), .ZN(n8414) );
  AOI22_X1 U1245 ( .A1(reg_mem[1304]), .A2(n3815), .B1(n8422), .B2(data_w[0]), 
        .ZN(n3814) );
  INV_X1 U1246 ( .A(n3816), .ZN(n8415) );
  AOI22_X1 U1247 ( .A1(reg_mem[1305]), .A2(n3815), .B1(n8422), .B2(data_w[1]), 
        .ZN(n3816) );
  INV_X1 U1248 ( .A(n3817), .ZN(n8416) );
  AOI22_X1 U1249 ( .A1(reg_mem[1306]), .A2(n3815), .B1(n8422), .B2(data_w[2]), 
        .ZN(n3817) );
  INV_X1 U1250 ( .A(n3818), .ZN(n8417) );
  AOI22_X1 U1251 ( .A1(reg_mem[1307]), .A2(n3815), .B1(n8422), .B2(data_w[3]), 
        .ZN(n3818) );
  INV_X1 U1252 ( .A(n3819), .ZN(n8418) );
  AOI22_X1 U1253 ( .A1(reg_mem[1308]), .A2(n3815), .B1(n8422), .B2(data_w[4]), 
        .ZN(n3819) );
  INV_X1 U1254 ( .A(n3820), .ZN(n8419) );
  AOI22_X1 U1255 ( .A1(reg_mem[1309]), .A2(n3815), .B1(n8422), .B2(data_w[5]), 
        .ZN(n3820) );
  INV_X1 U1256 ( .A(n3821), .ZN(n8420) );
  AOI22_X1 U1257 ( .A1(reg_mem[1310]), .A2(n3815), .B1(n8422), .B2(data_w[6]), 
        .ZN(n3821) );
  INV_X1 U1258 ( .A(n3822), .ZN(n8421) );
  AOI22_X1 U1259 ( .A1(reg_mem[1311]), .A2(n3815), .B1(n8422), .B2(data_w[7]), 
        .ZN(n3822) );
  INV_X1 U1260 ( .A(n3823), .ZN(n7117) );
  AOI22_X1 U1261 ( .A1(reg_mem[1312]), .A2(n3824), .B1(n7125), .B2(data_w[0]), 
        .ZN(n3823) );
  INV_X1 U1262 ( .A(n3825), .ZN(n7118) );
  AOI22_X1 U1263 ( .A1(reg_mem[1313]), .A2(n3824), .B1(n7125), .B2(data_w[1]), 
        .ZN(n3825) );
  INV_X1 U1264 ( .A(n3826), .ZN(n7119) );
  AOI22_X1 U1265 ( .A1(reg_mem[1314]), .A2(n3824), .B1(n7125), .B2(data_w[2]), 
        .ZN(n3826) );
  INV_X1 U1266 ( .A(n3827), .ZN(n7120) );
  AOI22_X1 U1267 ( .A1(reg_mem[1315]), .A2(n3824), .B1(n7125), .B2(data_w[3]), 
        .ZN(n3827) );
  INV_X1 U1268 ( .A(n3828), .ZN(n7121) );
  AOI22_X1 U1269 ( .A1(reg_mem[1316]), .A2(n3824), .B1(n7125), .B2(data_w[4]), 
        .ZN(n3828) );
  INV_X1 U1270 ( .A(n3829), .ZN(n7122) );
  AOI22_X1 U1271 ( .A1(reg_mem[1317]), .A2(n3824), .B1(n7125), .B2(data_w[5]), 
        .ZN(n3829) );
  INV_X1 U1272 ( .A(n3830), .ZN(n7123) );
  AOI22_X1 U1273 ( .A1(reg_mem[1318]), .A2(n3824), .B1(n7125), .B2(data_w[6]), 
        .ZN(n3830) );
  INV_X1 U1274 ( .A(n3831), .ZN(n7124) );
  AOI22_X1 U1275 ( .A1(reg_mem[1319]), .A2(n3824), .B1(n7125), .B2(data_w[7]), 
        .ZN(n3831) );
  INV_X1 U1276 ( .A(n3832), .ZN(n8846) );
  AOI22_X1 U1277 ( .A1(reg_mem[1320]), .A2(n3833), .B1(n8854), .B2(data_w[0]), 
        .ZN(n3832) );
  INV_X1 U1278 ( .A(n3834), .ZN(n8847) );
  AOI22_X1 U1279 ( .A1(reg_mem[1321]), .A2(n3833), .B1(n8854), .B2(data_w[1]), 
        .ZN(n3834) );
  INV_X1 U1280 ( .A(n3835), .ZN(n8848) );
  AOI22_X1 U1281 ( .A1(reg_mem[1322]), .A2(n3833), .B1(n8854), .B2(data_w[2]), 
        .ZN(n3835) );
  INV_X1 U1282 ( .A(n3836), .ZN(n8849) );
  AOI22_X1 U1283 ( .A1(reg_mem[1323]), .A2(n3833), .B1(n8854), .B2(data_w[3]), 
        .ZN(n3836) );
  INV_X1 U1284 ( .A(n3837), .ZN(n8850) );
  AOI22_X1 U1285 ( .A1(reg_mem[1324]), .A2(n3833), .B1(n8854), .B2(data_w[4]), 
        .ZN(n3837) );
  INV_X1 U1286 ( .A(n3838), .ZN(n8851) );
  AOI22_X1 U1287 ( .A1(reg_mem[1325]), .A2(n3833), .B1(n8854), .B2(data_w[5]), 
        .ZN(n3838) );
  INV_X1 U1288 ( .A(n3839), .ZN(n8852) );
  AOI22_X1 U1289 ( .A1(reg_mem[1326]), .A2(n3833), .B1(n8854), .B2(data_w[6]), 
        .ZN(n3839) );
  INV_X1 U1290 ( .A(n3840), .ZN(n8853) );
  AOI22_X1 U1291 ( .A1(reg_mem[1327]), .A2(n3833), .B1(n8854), .B2(data_w[7]), 
        .ZN(n3840) );
  INV_X1 U1292 ( .A(n3841), .ZN(n7693) );
  AOI22_X1 U1293 ( .A1(reg_mem[1328]), .A2(n3842), .B1(n7701), .B2(data_w[0]), 
        .ZN(n3841) );
  INV_X1 U1294 ( .A(n3843), .ZN(n7694) );
  AOI22_X1 U1295 ( .A1(reg_mem[1329]), .A2(n3842), .B1(n7701), .B2(data_w[1]), 
        .ZN(n3843) );
  INV_X1 U1296 ( .A(n3844), .ZN(n7695) );
  AOI22_X1 U1297 ( .A1(reg_mem[1330]), .A2(n3842), .B1(n7701), .B2(data_w[2]), 
        .ZN(n3844) );
  INV_X1 U1298 ( .A(n3845), .ZN(n7696) );
  AOI22_X1 U1299 ( .A1(reg_mem[1331]), .A2(n3842), .B1(n7701), .B2(data_w[3]), 
        .ZN(n3845) );
  INV_X1 U1300 ( .A(n3846), .ZN(n7697) );
  AOI22_X1 U1301 ( .A1(reg_mem[1332]), .A2(n3842), .B1(n7701), .B2(data_w[4]), 
        .ZN(n3846) );
  INV_X1 U1302 ( .A(n3847), .ZN(n7698) );
  AOI22_X1 U1303 ( .A1(reg_mem[1333]), .A2(n3842), .B1(n7701), .B2(data_w[5]), 
        .ZN(n3847) );
  INV_X1 U1304 ( .A(n3848), .ZN(n7699) );
  AOI22_X1 U1305 ( .A1(reg_mem[1334]), .A2(n3842), .B1(n7701), .B2(data_w[6]), 
        .ZN(n3848) );
  INV_X1 U1306 ( .A(n3849), .ZN(n7700) );
  AOI22_X1 U1307 ( .A1(reg_mem[1335]), .A2(n3842), .B1(n7701), .B2(data_w[7]), 
        .ZN(n3849) );
  INV_X1 U1308 ( .A(n3850), .ZN(n8270) );
  AOI22_X1 U1309 ( .A1(reg_mem[1336]), .A2(n3851), .B1(n8278), .B2(data_w[0]), 
        .ZN(n3850) );
  INV_X1 U1310 ( .A(n3852), .ZN(n8271) );
  AOI22_X1 U1311 ( .A1(reg_mem[1337]), .A2(n3851), .B1(n8278), .B2(data_w[1]), 
        .ZN(n3852) );
  INV_X1 U1312 ( .A(n3853), .ZN(n8272) );
  AOI22_X1 U1313 ( .A1(reg_mem[1338]), .A2(n3851), .B1(n8278), .B2(data_w[2]), 
        .ZN(n3853) );
  INV_X1 U1314 ( .A(n3854), .ZN(n8273) );
  AOI22_X1 U1315 ( .A1(reg_mem[1339]), .A2(n3851), .B1(n8278), .B2(data_w[3]), 
        .ZN(n3854) );
  INV_X1 U1316 ( .A(n3855), .ZN(n8274) );
  AOI22_X1 U1317 ( .A1(reg_mem[1340]), .A2(n3851), .B1(n8278), .B2(data_w[4]), 
        .ZN(n3855) );
  INV_X1 U1318 ( .A(n3856), .ZN(n8275) );
  AOI22_X1 U1319 ( .A1(reg_mem[1341]), .A2(n3851), .B1(n8278), .B2(data_w[5]), 
        .ZN(n3856) );
  INV_X1 U1320 ( .A(n3857), .ZN(n8276) );
  AOI22_X1 U1321 ( .A1(reg_mem[1342]), .A2(n3851), .B1(n8278), .B2(data_w[6]), 
        .ZN(n3857) );
  INV_X1 U1322 ( .A(n3858), .ZN(n8277) );
  AOI22_X1 U1323 ( .A1(reg_mem[1343]), .A2(n3851), .B1(n8278), .B2(data_w[7]), 
        .ZN(n3858) );
  INV_X1 U1324 ( .A(n3859), .ZN(n6973) );
  AOI22_X1 U1325 ( .A1(reg_mem[1344]), .A2(n3860), .B1(n6981), .B2(data_w[0]), 
        .ZN(n3859) );
  INV_X1 U1326 ( .A(n3861), .ZN(n6974) );
  AOI22_X1 U1327 ( .A1(reg_mem[1345]), .A2(n3860), .B1(n6981), .B2(data_w[1]), 
        .ZN(n3861) );
  INV_X1 U1328 ( .A(n3862), .ZN(n6975) );
  AOI22_X1 U1329 ( .A1(reg_mem[1346]), .A2(n3860), .B1(n6981), .B2(data_w[2]), 
        .ZN(n3862) );
  INV_X1 U1330 ( .A(n3863), .ZN(n6976) );
  AOI22_X1 U1331 ( .A1(reg_mem[1347]), .A2(n3860), .B1(n6981), .B2(data_w[3]), 
        .ZN(n3863) );
  INV_X1 U1332 ( .A(n3864), .ZN(n6977) );
  AOI22_X1 U1333 ( .A1(reg_mem[1348]), .A2(n3860), .B1(n6981), .B2(data_w[4]), 
        .ZN(n3864) );
  INV_X1 U1334 ( .A(n3865), .ZN(n6978) );
  AOI22_X1 U1335 ( .A1(reg_mem[1349]), .A2(n3860), .B1(n6981), .B2(data_w[5]), 
        .ZN(n3865) );
  INV_X1 U1336 ( .A(n3866), .ZN(n6979) );
  AOI22_X1 U1337 ( .A1(reg_mem[1350]), .A2(n3860), .B1(n6981), .B2(data_w[6]), 
        .ZN(n3866) );
  INV_X1 U1338 ( .A(n3867), .ZN(n6980) );
  AOI22_X1 U1339 ( .A1(reg_mem[1351]), .A2(n3860), .B1(n6981), .B2(data_w[7]), 
        .ZN(n3867) );
  INV_X1 U1340 ( .A(n3868), .ZN(n8702) );
  AOI22_X1 U1341 ( .A1(reg_mem[1352]), .A2(n3869), .B1(n8710), .B2(data_w[0]), 
        .ZN(n3868) );
  INV_X1 U1342 ( .A(n3870), .ZN(n8703) );
  AOI22_X1 U1343 ( .A1(reg_mem[1353]), .A2(n3869), .B1(n8710), .B2(data_w[1]), 
        .ZN(n3870) );
  INV_X1 U1344 ( .A(n3871), .ZN(n8704) );
  AOI22_X1 U1345 ( .A1(reg_mem[1354]), .A2(n3869), .B1(n8710), .B2(data_w[2]), 
        .ZN(n3871) );
  INV_X1 U1346 ( .A(n3872), .ZN(n8705) );
  AOI22_X1 U1347 ( .A1(reg_mem[1355]), .A2(n3869), .B1(n8710), .B2(data_w[3]), 
        .ZN(n3872) );
  INV_X1 U1348 ( .A(n3873), .ZN(n8706) );
  AOI22_X1 U1349 ( .A1(reg_mem[1356]), .A2(n3869), .B1(n8710), .B2(data_w[4]), 
        .ZN(n3873) );
  INV_X1 U1350 ( .A(n3874), .ZN(n8707) );
  AOI22_X1 U1351 ( .A1(reg_mem[1357]), .A2(n3869), .B1(n8710), .B2(data_w[5]), 
        .ZN(n3874) );
  INV_X1 U1352 ( .A(n3875), .ZN(n8708) );
  AOI22_X1 U1353 ( .A1(reg_mem[1358]), .A2(n3869), .B1(n8710), .B2(data_w[6]), 
        .ZN(n3875) );
  INV_X1 U1354 ( .A(n3876), .ZN(n8709) );
  AOI22_X1 U1355 ( .A1(reg_mem[1359]), .A2(n3869), .B1(n8710), .B2(data_w[7]), 
        .ZN(n3876) );
  INV_X1 U1356 ( .A(n3877), .ZN(n7549) );
  AOI22_X1 U1357 ( .A1(reg_mem[1360]), .A2(n3878), .B1(n7557), .B2(data_w[0]), 
        .ZN(n3877) );
  INV_X1 U1358 ( .A(n3879), .ZN(n7550) );
  AOI22_X1 U1359 ( .A1(reg_mem[1361]), .A2(n3878), .B1(n7557), .B2(data_w[1]), 
        .ZN(n3879) );
  INV_X1 U1360 ( .A(n3880), .ZN(n7551) );
  AOI22_X1 U1361 ( .A1(reg_mem[1362]), .A2(n3878), .B1(n7557), .B2(data_w[2]), 
        .ZN(n3880) );
  INV_X1 U1362 ( .A(n3881), .ZN(n7552) );
  AOI22_X1 U1363 ( .A1(reg_mem[1363]), .A2(n3878), .B1(n7557), .B2(data_w[3]), 
        .ZN(n3881) );
  INV_X1 U1364 ( .A(n3882), .ZN(n7553) );
  AOI22_X1 U1365 ( .A1(reg_mem[1364]), .A2(n3878), .B1(n7557), .B2(data_w[4]), 
        .ZN(n3882) );
  INV_X1 U1366 ( .A(n3883), .ZN(n7554) );
  AOI22_X1 U1367 ( .A1(reg_mem[1365]), .A2(n3878), .B1(n7557), .B2(data_w[5]), 
        .ZN(n3883) );
  INV_X1 U1368 ( .A(n3884), .ZN(n7555) );
  AOI22_X1 U1369 ( .A1(reg_mem[1366]), .A2(n3878), .B1(n7557), .B2(data_w[6]), 
        .ZN(n3884) );
  INV_X1 U1370 ( .A(n3885), .ZN(n7556) );
  AOI22_X1 U1371 ( .A1(reg_mem[1367]), .A2(n3878), .B1(n7557), .B2(data_w[7]), 
        .ZN(n3885) );
  INV_X1 U1372 ( .A(n3886), .ZN(n8126) );
  AOI22_X1 U1373 ( .A1(reg_mem[1368]), .A2(n3887), .B1(n8134), .B2(data_w[0]), 
        .ZN(n3886) );
  INV_X1 U1374 ( .A(n3888), .ZN(n8127) );
  AOI22_X1 U1375 ( .A1(reg_mem[1369]), .A2(n3887), .B1(n8134), .B2(data_w[1]), 
        .ZN(n3888) );
  INV_X1 U1376 ( .A(n3889), .ZN(n8128) );
  AOI22_X1 U1377 ( .A1(reg_mem[1370]), .A2(n3887), .B1(n8134), .B2(data_w[2]), 
        .ZN(n3889) );
  INV_X1 U1378 ( .A(n3890), .ZN(n8129) );
  AOI22_X1 U1379 ( .A1(reg_mem[1371]), .A2(n3887), .B1(n8134), .B2(data_w[3]), 
        .ZN(n3890) );
  INV_X1 U1380 ( .A(n3891), .ZN(n8130) );
  AOI22_X1 U1381 ( .A1(reg_mem[1372]), .A2(n3887), .B1(n8134), .B2(data_w[4]), 
        .ZN(n3891) );
  INV_X1 U1382 ( .A(n3892), .ZN(n8131) );
  AOI22_X1 U1383 ( .A1(reg_mem[1373]), .A2(n3887), .B1(n8134), .B2(data_w[5]), 
        .ZN(n3892) );
  INV_X1 U1384 ( .A(n3893), .ZN(n8132) );
  AOI22_X1 U1385 ( .A1(reg_mem[1374]), .A2(n3887), .B1(n8134), .B2(data_w[6]), 
        .ZN(n3893) );
  INV_X1 U1386 ( .A(n3894), .ZN(n8133) );
  AOI22_X1 U1387 ( .A1(reg_mem[1375]), .A2(n3887), .B1(n8134), .B2(data_w[7]), 
        .ZN(n3894) );
  INV_X1 U1388 ( .A(n2324), .ZN(n9080) );
  AOI22_X1 U1389 ( .A1(reg_mem[8]), .A2(n2325), .B1(n9088), .B2(data_w[0]), 
        .ZN(n2324) );
  INV_X1 U1390 ( .A(n2326), .ZN(n9081) );
  AOI22_X1 U1391 ( .A1(reg_mem[9]), .A2(n2325), .B1(n9088), .B2(data_w[1]), 
        .ZN(n2326) );
  INV_X1 U1392 ( .A(n2327), .ZN(n9082) );
  AOI22_X1 U1393 ( .A1(reg_mem[10]), .A2(n2325), .B1(n9088), .B2(data_w[2]), 
        .ZN(n2327) );
  INV_X1 U1394 ( .A(n2328), .ZN(n9083) );
  AOI22_X1 U1395 ( .A1(reg_mem[11]), .A2(n2325), .B1(n9088), .B2(data_w[3]), 
        .ZN(n2328) );
  INV_X1 U1396 ( .A(n2329), .ZN(n9084) );
  AOI22_X1 U1397 ( .A1(reg_mem[12]), .A2(n2325), .B1(n9088), .B2(data_w[4]), 
        .ZN(n2329) );
  INV_X1 U1398 ( .A(n2330), .ZN(n9085) );
  AOI22_X1 U1399 ( .A1(reg_mem[13]), .A2(n2325), .B1(n9088), .B2(data_w[5]), 
        .ZN(n2330) );
  INV_X1 U1400 ( .A(n2331), .ZN(n9086) );
  AOI22_X1 U1401 ( .A1(reg_mem[14]), .A2(n2325), .B1(n9088), .B2(data_w[6]), 
        .ZN(n2331) );
  INV_X1 U1402 ( .A(n2332), .ZN(n9087) );
  AOI22_X1 U1403 ( .A1(reg_mem[15]), .A2(n2325), .B1(n9088), .B2(data_w[7]), 
        .ZN(n2332) );
  INV_X1 U1404 ( .A(n2334), .ZN(n7927) );
  AOI22_X1 U1405 ( .A1(reg_mem[16]), .A2(n2335), .B1(n7935), .B2(data_w[0]), 
        .ZN(n2334) );
  INV_X1 U1406 ( .A(n2336), .ZN(n7928) );
  AOI22_X1 U1407 ( .A1(reg_mem[17]), .A2(n2335), .B1(n7935), .B2(data_w[1]), 
        .ZN(n2336) );
  INV_X1 U1408 ( .A(n2337), .ZN(n7929) );
  AOI22_X1 U1409 ( .A1(reg_mem[18]), .A2(n2335), .B1(n7935), .B2(data_w[2]), 
        .ZN(n2337) );
  INV_X1 U1410 ( .A(n2338), .ZN(n7930) );
  AOI22_X1 U1411 ( .A1(reg_mem[19]), .A2(n2335), .B1(n7935), .B2(data_w[3]), 
        .ZN(n2338) );
  INV_X1 U1412 ( .A(n2339), .ZN(n7931) );
  AOI22_X1 U1413 ( .A1(reg_mem[20]), .A2(n2335), .B1(n7935), .B2(data_w[4]), 
        .ZN(n2339) );
  INV_X1 U1414 ( .A(n2340), .ZN(n7932) );
  AOI22_X1 U1415 ( .A1(reg_mem[21]), .A2(n2335), .B1(n7935), .B2(data_w[5]), 
        .ZN(n2340) );
  INV_X1 U1416 ( .A(n2341), .ZN(n7933) );
  AOI22_X1 U1417 ( .A1(reg_mem[22]), .A2(n2335), .B1(n7935), .B2(data_w[6]), 
        .ZN(n2341) );
  INV_X1 U1418 ( .A(n2342), .ZN(n7934) );
  AOI22_X1 U1419 ( .A1(reg_mem[23]), .A2(n2335), .B1(n7935), .B2(data_w[7]), 
        .ZN(n2342) );
  INV_X1 U1420 ( .A(n2344), .ZN(n8504) );
  AOI22_X1 U1421 ( .A1(reg_mem[24]), .A2(n2345), .B1(n8512), .B2(data_w[0]), 
        .ZN(n2344) );
  INV_X1 U1422 ( .A(n2346), .ZN(n8505) );
  AOI22_X1 U1423 ( .A1(reg_mem[25]), .A2(n2345), .B1(n8512), .B2(data_w[1]), 
        .ZN(n2346) );
  INV_X1 U1424 ( .A(n2347), .ZN(n8506) );
  AOI22_X1 U1425 ( .A1(reg_mem[26]), .A2(n2345), .B1(n8512), .B2(data_w[2]), 
        .ZN(n2347) );
  INV_X1 U1426 ( .A(n2348), .ZN(n8507) );
  AOI22_X1 U1427 ( .A1(reg_mem[27]), .A2(n2345), .B1(n8512), .B2(data_w[3]), 
        .ZN(n2348) );
  INV_X1 U1428 ( .A(n2349), .ZN(n8508) );
  AOI22_X1 U1429 ( .A1(reg_mem[28]), .A2(n2345), .B1(n8512), .B2(data_w[4]), 
        .ZN(n2349) );
  INV_X1 U1430 ( .A(n2350), .ZN(n8509) );
  AOI22_X1 U1431 ( .A1(reg_mem[29]), .A2(n2345), .B1(n8512), .B2(data_w[5]), 
        .ZN(n2350) );
  INV_X1 U1432 ( .A(n2351), .ZN(n8510) );
  AOI22_X1 U1433 ( .A1(reg_mem[30]), .A2(n2345), .B1(n8512), .B2(data_w[6]), 
        .ZN(n2351) );
  INV_X1 U1434 ( .A(n2352), .ZN(n8511) );
  AOI22_X1 U1435 ( .A1(reg_mem[31]), .A2(n2345), .B1(n8512), .B2(data_w[7]), 
        .ZN(n2352) );
  INV_X1 U1436 ( .A(n2805), .ZN(n7180) );
  AOI22_X1 U1437 ( .A1(reg_mem[416]), .A2(n2806), .B1(n7188), .B2(data_w[0]), 
        .ZN(n2805) );
  INV_X1 U1438 ( .A(n2807), .ZN(n7181) );
  AOI22_X1 U1439 ( .A1(reg_mem[417]), .A2(n2806), .B1(n7188), .B2(data_w[1]), 
        .ZN(n2807) );
  INV_X1 U1440 ( .A(n2808), .ZN(n7182) );
  AOI22_X1 U1441 ( .A1(reg_mem[418]), .A2(n2806), .B1(n7188), .B2(data_w[2]), 
        .ZN(n2808) );
  INV_X1 U1442 ( .A(n2809), .ZN(n7183) );
  AOI22_X1 U1443 ( .A1(reg_mem[419]), .A2(n2806), .B1(n7188), .B2(data_w[3]), 
        .ZN(n2809) );
  INV_X1 U1444 ( .A(n2810), .ZN(n7184) );
  AOI22_X1 U1445 ( .A1(reg_mem[420]), .A2(n2806), .B1(n7188), .B2(data_w[4]), 
        .ZN(n2810) );
  INV_X1 U1446 ( .A(n2811), .ZN(n7185) );
  AOI22_X1 U1447 ( .A1(reg_mem[421]), .A2(n2806), .B1(n7188), .B2(data_w[5]), 
        .ZN(n2811) );
  INV_X1 U1448 ( .A(n2812), .ZN(n7186) );
  AOI22_X1 U1449 ( .A1(reg_mem[422]), .A2(n2806), .B1(n7188), .B2(data_w[6]), 
        .ZN(n2812) );
  INV_X1 U1450 ( .A(n2813), .ZN(n7187) );
  AOI22_X1 U1451 ( .A1(reg_mem[423]), .A2(n2806), .B1(n7188), .B2(data_w[7]), 
        .ZN(n2813) );
  INV_X1 U1452 ( .A(n2814), .ZN(n8909) );
  AOI22_X1 U1453 ( .A1(reg_mem[424]), .A2(n2815), .B1(n8917), .B2(data_w[0]), 
        .ZN(n2814) );
  INV_X1 U1454 ( .A(n2816), .ZN(n8910) );
  AOI22_X1 U1455 ( .A1(reg_mem[425]), .A2(n2815), .B1(n8917), .B2(data_w[1]), 
        .ZN(n2816) );
  INV_X1 U1456 ( .A(n2817), .ZN(n8911) );
  AOI22_X1 U1457 ( .A1(reg_mem[426]), .A2(n2815), .B1(n8917), .B2(data_w[2]), 
        .ZN(n2817) );
  INV_X1 U1458 ( .A(n2818), .ZN(n8912) );
  AOI22_X1 U1459 ( .A1(reg_mem[427]), .A2(n2815), .B1(n8917), .B2(data_w[3]), 
        .ZN(n2818) );
  INV_X1 U1460 ( .A(n2819), .ZN(n8913) );
  AOI22_X1 U1461 ( .A1(reg_mem[428]), .A2(n2815), .B1(n8917), .B2(data_w[4]), 
        .ZN(n2819) );
  INV_X1 U1462 ( .A(n2820), .ZN(n8914) );
  AOI22_X1 U1463 ( .A1(reg_mem[429]), .A2(n2815), .B1(n8917), .B2(data_w[5]), 
        .ZN(n2820) );
  INV_X1 U1464 ( .A(n2821), .ZN(n8915) );
  AOI22_X1 U1465 ( .A1(reg_mem[430]), .A2(n2815), .B1(n8917), .B2(data_w[6]), 
        .ZN(n2821) );
  INV_X1 U1466 ( .A(n2822), .ZN(n8916) );
  AOI22_X1 U1467 ( .A1(reg_mem[431]), .A2(n2815), .B1(n8917), .B2(data_w[7]), 
        .ZN(n2822) );
  INV_X1 U1468 ( .A(n2823), .ZN(n7756) );
  AOI22_X1 U1469 ( .A1(reg_mem[432]), .A2(n2824), .B1(n7764), .B2(data_w[0]), 
        .ZN(n2823) );
  INV_X1 U1470 ( .A(n2825), .ZN(n7757) );
  AOI22_X1 U1471 ( .A1(reg_mem[433]), .A2(n2824), .B1(n7764), .B2(data_w[1]), 
        .ZN(n2825) );
  INV_X1 U1472 ( .A(n2826), .ZN(n7758) );
  AOI22_X1 U1473 ( .A1(reg_mem[434]), .A2(n2824), .B1(n7764), .B2(data_w[2]), 
        .ZN(n2826) );
  INV_X1 U1474 ( .A(n2827), .ZN(n7759) );
  AOI22_X1 U1475 ( .A1(reg_mem[435]), .A2(n2824), .B1(n7764), .B2(data_w[3]), 
        .ZN(n2827) );
  INV_X1 U1476 ( .A(n2828), .ZN(n7760) );
  AOI22_X1 U1477 ( .A1(reg_mem[436]), .A2(n2824), .B1(n7764), .B2(data_w[4]), 
        .ZN(n2828) );
  INV_X1 U1478 ( .A(n2829), .ZN(n7761) );
  AOI22_X1 U1479 ( .A1(reg_mem[437]), .A2(n2824), .B1(n7764), .B2(data_w[5]), 
        .ZN(n2829) );
  INV_X1 U1480 ( .A(n2830), .ZN(n7762) );
  AOI22_X1 U1481 ( .A1(reg_mem[438]), .A2(n2824), .B1(n7764), .B2(data_w[6]), 
        .ZN(n2830) );
  INV_X1 U1482 ( .A(n2831), .ZN(n7763) );
  AOI22_X1 U1483 ( .A1(reg_mem[439]), .A2(n2824), .B1(n7764), .B2(data_w[7]), 
        .ZN(n2831) );
  INV_X1 U1484 ( .A(n2832), .ZN(n8333) );
  AOI22_X1 U1485 ( .A1(reg_mem[440]), .A2(n2833), .B1(n8341), .B2(data_w[0]), 
        .ZN(n2832) );
  INV_X1 U1486 ( .A(n2834), .ZN(n8334) );
  AOI22_X1 U1487 ( .A1(reg_mem[441]), .A2(n2833), .B1(n8341), .B2(data_w[1]), 
        .ZN(n2834) );
  INV_X1 U1488 ( .A(n2835), .ZN(n8335) );
  AOI22_X1 U1489 ( .A1(reg_mem[442]), .A2(n2833), .B1(n8341), .B2(data_w[2]), 
        .ZN(n2835) );
  INV_X1 U1490 ( .A(n2836), .ZN(n8336) );
  AOI22_X1 U1491 ( .A1(reg_mem[443]), .A2(n2833), .B1(n8341), .B2(data_w[3]), 
        .ZN(n2836) );
  INV_X1 U1492 ( .A(n2837), .ZN(n8337) );
  AOI22_X1 U1493 ( .A1(reg_mem[444]), .A2(n2833), .B1(n8341), .B2(data_w[4]), 
        .ZN(n2837) );
  INV_X1 U1494 ( .A(n2838), .ZN(n8338) );
  AOI22_X1 U1495 ( .A1(reg_mem[445]), .A2(n2833), .B1(n8341), .B2(data_w[5]), 
        .ZN(n2838) );
  INV_X1 U1496 ( .A(n2839), .ZN(n8339) );
  AOI22_X1 U1497 ( .A1(reg_mem[446]), .A2(n2833), .B1(n8341), .B2(data_w[6]), 
        .ZN(n2839) );
  INV_X1 U1498 ( .A(n2840), .ZN(n8340) );
  AOI22_X1 U1499 ( .A1(reg_mem[447]), .A2(n2833), .B1(n8341), .B2(data_w[7]), 
        .ZN(n2840) );
  INV_X1 U1500 ( .A(n2841), .ZN(n7036) );
  AOI22_X1 U1501 ( .A1(reg_mem[448]), .A2(n2842), .B1(n7044), .B2(data_w[0]), 
        .ZN(n2841) );
  INV_X1 U1502 ( .A(n2843), .ZN(n7037) );
  AOI22_X1 U1503 ( .A1(reg_mem[449]), .A2(n2842), .B1(n7044), .B2(data_w[1]), 
        .ZN(n2843) );
  INV_X1 U1504 ( .A(n2844), .ZN(n7038) );
  AOI22_X1 U1505 ( .A1(reg_mem[450]), .A2(n2842), .B1(n7044), .B2(data_w[2]), 
        .ZN(n2844) );
  INV_X1 U1506 ( .A(n2845), .ZN(n7039) );
  AOI22_X1 U1507 ( .A1(reg_mem[451]), .A2(n2842), .B1(n7044), .B2(data_w[3]), 
        .ZN(n2845) );
  INV_X1 U1508 ( .A(n2846), .ZN(n7040) );
  AOI22_X1 U1509 ( .A1(reg_mem[452]), .A2(n2842), .B1(n7044), .B2(data_w[4]), 
        .ZN(n2846) );
  INV_X1 U1510 ( .A(n2847), .ZN(n7041) );
  AOI22_X1 U1511 ( .A1(reg_mem[453]), .A2(n2842), .B1(n7044), .B2(data_w[5]), 
        .ZN(n2847) );
  INV_X1 U1512 ( .A(n2848), .ZN(n7042) );
  AOI22_X1 U1513 ( .A1(reg_mem[454]), .A2(n2842), .B1(n7044), .B2(data_w[6]), 
        .ZN(n2848) );
  INV_X1 U1514 ( .A(n2849), .ZN(n7043) );
  AOI22_X1 U1515 ( .A1(reg_mem[455]), .A2(n2842), .B1(n7044), .B2(data_w[7]), 
        .ZN(n2849) );
  INV_X1 U1516 ( .A(n2850), .ZN(n8765) );
  AOI22_X1 U1517 ( .A1(reg_mem[456]), .A2(n2851), .B1(n8773), .B2(data_w[0]), 
        .ZN(n2850) );
  INV_X1 U1518 ( .A(n2852), .ZN(n8766) );
  AOI22_X1 U1519 ( .A1(reg_mem[457]), .A2(n2851), .B1(n8773), .B2(data_w[1]), 
        .ZN(n2852) );
  INV_X1 U1520 ( .A(n2853), .ZN(n8767) );
  AOI22_X1 U1521 ( .A1(reg_mem[458]), .A2(n2851), .B1(n8773), .B2(data_w[2]), 
        .ZN(n2853) );
  INV_X1 U1522 ( .A(n2854), .ZN(n8768) );
  AOI22_X1 U1523 ( .A1(reg_mem[459]), .A2(n2851), .B1(n8773), .B2(data_w[3]), 
        .ZN(n2854) );
  INV_X1 U1524 ( .A(n2855), .ZN(n8769) );
  AOI22_X1 U1525 ( .A1(reg_mem[460]), .A2(n2851), .B1(n8773), .B2(data_w[4]), 
        .ZN(n2855) );
  INV_X1 U1526 ( .A(n2856), .ZN(n8770) );
  AOI22_X1 U1527 ( .A1(reg_mem[461]), .A2(n2851), .B1(n8773), .B2(data_w[5]), 
        .ZN(n2856) );
  INV_X1 U1528 ( .A(n2857), .ZN(n8771) );
  AOI22_X1 U1529 ( .A1(reg_mem[462]), .A2(n2851), .B1(n8773), .B2(data_w[6]), 
        .ZN(n2857) );
  INV_X1 U1530 ( .A(n2858), .ZN(n8772) );
  AOI22_X1 U1531 ( .A1(reg_mem[463]), .A2(n2851), .B1(n8773), .B2(data_w[7]), 
        .ZN(n2858) );
  INV_X1 U1532 ( .A(n2859), .ZN(n7612) );
  AOI22_X1 U1533 ( .A1(reg_mem[464]), .A2(n2860), .B1(n7620), .B2(data_w[0]), 
        .ZN(n2859) );
  INV_X1 U1534 ( .A(n2861), .ZN(n7613) );
  AOI22_X1 U1535 ( .A1(reg_mem[465]), .A2(n2860), .B1(n7620), .B2(data_w[1]), 
        .ZN(n2861) );
  INV_X1 U1536 ( .A(n2862), .ZN(n7614) );
  AOI22_X1 U1537 ( .A1(reg_mem[466]), .A2(n2860), .B1(n7620), .B2(data_w[2]), 
        .ZN(n2862) );
  INV_X1 U1538 ( .A(n2863), .ZN(n7615) );
  AOI22_X1 U1539 ( .A1(reg_mem[467]), .A2(n2860), .B1(n7620), .B2(data_w[3]), 
        .ZN(n2863) );
  INV_X1 U1540 ( .A(n2864), .ZN(n7616) );
  AOI22_X1 U1541 ( .A1(reg_mem[468]), .A2(n2860), .B1(n7620), .B2(data_w[4]), 
        .ZN(n2864) );
  INV_X1 U1542 ( .A(n2865), .ZN(n7617) );
  AOI22_X1 U1543 ( .A1(reg_mem[469]), .A2(n2860), .B1(n7620), .B2(data_w[5]), 
        .ZN(n2865) );
  INV_X1 U1544 ( .A(n2866), .ZN(n7618) );
  AOI22_X1 U1545 ( .A1(reg_mem[470]), .A2(n2860), .B1(n7620), .B2(data_w[6]), 
        .ZN(n2866) );
  INV_X1 U1546 ( .A(n2867), .ZN(n7619) );
  AOI22_X1 U1547 ( .A1(reg_mem[471]), .A2(n2860), .B1(n7620), .B2(data_w[7]), 
        .ZN(n2867) );
  INV_X1 U1548 ( .A(n2868), .ZN(n8189) );
  AOI22_X1 U1549 ( .A1(reg_mem[472]), .A2(n2869), .B1(n8197), .B2(data_w[0]), 
        .ZN(n2868) );
  INV_X1 U1550 ( .A(n2870), .ZN(n8190) );
  AOI22_X1 U1551 ( .A1(reg_mem[473]), .A2(n2869), .B1(n8197), .B2(data_w[1]), 
        .ZN(n2870) );
  INV_X1 U1552 ( .A(n2871), .ZN(n8191) );
  AOI22_X1 U1553 ( .A1(reg_mem[474]), .A2(n2869), .B1(n8197), .B2(data_w[2]), 
        .ZN(n2871) );
  INV_X1 U1554 ( .A(n2872), .ZN(n8192) );
  AOI22_X1 U1555 ( .A1(reg_mem[475]), .A2(n2869), .B1(n8197), .B2(data_w[3]), 
        .ZN(n2872) );
  INV_X1 U1556 ( .A(n2873), .ZN(n8193) );
  AOI22_X1 U1557 ( .A1(reg_mem[476]), .A2(n2869), .B1(n8197), .B2(data_w[4]), 
        .ZN(n2873) );
  INV_X1 U1558 ( .A(n2874), .ZN(n8194) );
  AOI22_X1 U1559 ( .A1(reg_mem[477]), .A2(n2869), .B1(n8197), .B2(data_w[5]), 
        .ZN(n2874) );
  INV_X1 U1560 ( .A(n2875), .ZN(n8195) );
  AOI22_X1 U1561 ( .A1(reg_mem[478]), .A2(n2869), .B1(n8197), .B2(data_w[6]), 
        .ZN(n2875) );
  INV_X1 U1562 ( .A(n2876), .ZN(n8196) );
  AOI22_X1 U1563 ( .A1(reg_mem[479]), .A2(n2869), .B1(n8197), .B2(data_w[7]), 
        .ZN(n2876) );
  INV_X1 U1564 ( .A(n2877), .ZN(n6892) );
  AOI22_X1 U1565 ( .A1(reg_mem[480]), .A2(n2878), .B1(n6900), .B2(data_w[0]), 
        .ZN(n2877) );
  INV_X1 U1566 ( .A(n2879), .ZN(n6893) );
  AOI22_X1 U1567 ( .A1(reg_mem[481]), .A2(n2878), .B1(n6900), .B2(data_w[1]), 
        .ZN(n2879) );
  INV_X1 U1568 ( .A(n2880), .ZN(n6894) );
  AOI22_X1 U1569 ( .A1(reg_mem[482]), .A2(n2878), .B1(n6900), .B2(data_w[2]), 
        .ZN(n2880) );
  INV_X1 U1570 ( .A(n2881), .ZN(n6895) );
  AOI22_X1 U1571 ( .A1(reg_mem[483]), .A2(n2878), .B1(n6900), .B2(data_w[3]), 
        .ZN(n2881) );
  INV_X1 U1572 ( .A(n2882), .ZN(n6896) );
  AOI22_X1 U1573 ( .A1(reg_mem[484]), .A2(n2878), .B1(n6900), .B2(data_w[4]), 
        .ZN(n2882) );
  INV_X1 U1574 ( .A(n2883), .ZN(n6897) );
  AOI22_X1 U1575 ( .A1(reg_mem[485]), .A2(n2878), .B1(n6900), .B2(data_w[5]), 
        .ZN(n2883) );
  INV_X1 U1576 ( .A(n2884), .ZN(n6898) );
  AOI22_X1 U1577 ( .A1(reg_mem[486]), .A2(n2878), .B1(n6900), .B2(data_w[6]), 
        .ZN(n2884) );
  INV_X1 U1578 ( .A(n2885), .ZN(n6899) );
  AOI22_X1 U1579 ( .A1(reg_mem[487]), .A2(n2878), .B1(n6900), .B2(data_w[7]), 
        .ZN(n2885) );
  INV_X1 U1580 ( .A(n2886), .ZN(n8621) );
  AOI22_X1 U1581 ( .A1(reg_mem[488]), .A2(n2887), .B1(n8629), .B2(data_w[0]), 
        .ZN(n2886) );
  INV_X1 U1582 ( .A(n2888), .ZN(n8622) );
  AOI22_X1 U1583 ( .A1(reg_mem[489]), .A2(n2887), .B1(n8629), .B2(data_w[1]), 
        .ZN(n2888) );
  INV_X1 U1584 ( .A(n2889), .ZN(n8623) );
  AOI22_X1 U1585 ( .A1(reg_mem[490]), .A2(n2887), .B1(n8629), .B2(data_w[2]), 
        .ZN(n2889) );
  INV_X1 U1586 ( .A(n2890), .ZN(n8624) );
  AOI22_X1 U1587 ( .A1(reg_mem[491]), .A2(n2887), .B1(n8629), .B2(data_w[3]), 
        .ZN(n2890) );
  INV_X1 U1588 ( .A(n2891), .ZN(n8625) );
  AOI22_X1 U1589 ( .A1(reg_mem[492]), .A2(n2887), .B1(n8629), .B2(data_w[4]), 
        .ZN(n2891) );
  INV_X1 U1590 ( .A(n2892), .ZN(n8626) );
  AOI22_X1 U1591 ( .A1(reg_mem[493]), .A2(n2887), .B1(n8629), .B2(data_w[5]), 
        .ZN(n2892) );
  INV_X1 U1592 ( .A(n2893), .ZN(n8627) );
  AOI22_X1 U1593 ( .A1(reg_mem[494]), .A2(n2887), .B1(n8629), .B2(data_w[6]), 
        .ZN(n2893) );
  INV_X1 U1594 ( .A(n2894), .ZN(n8628) );
  AOI22_X1 U1595 ( .A1(reg_mem[495]), .A2(n2887), .B1(n8629), .B2(data_w[7]), 
        .ZN(n2894) );
  INV_X1 U1596 ( .A(n2895), .ZN(n7468) );
  AOI22_X1 U1597 ( .A1(reg_mem[496]), .A2(n2896), .B1(n7476), .B2(data_w[0]), 
        .ZN(n2895) );
  INV_X1 U1598 ( .A(n2897), .ZN(n7469) );
  AOI22_X1 U1599 ( .A1(reg_mem[497]), .A2(n2896), .B1(n7476), .B2(data_w[1]), 
        .ZN(n2897) );
  INV_X1 U1600 ( .A(n2898), .ZN(n7470) );
  AOI22_X1 U1601 ( .A1(reg_mem[498]), .A2(n2896), .B1(n7476), .B2(data_w[2]), 
        .ZN(n2898) );
  INV_X1 U1602 ( .A(n2899), .ZN(n7471) );
  AOI22_X1 U1603 ( .A1(reg_mem[499]), .A2(n2896), .B1(n7476), .B2(data_w[3]), 
        .ZN(n2899) );
  INV_X1 U1604 ( .A(n2900), .ZN(n7472) );
  AOI22_X1 U1605 ( .A1(reg_mem[500]), .A2(n2896), .B1(n7476), .B2(data_w[4]), 
        .ZN(n2900) );
  INV_X1 U1606 ( .A(n2901), .ZN(n7473) );
  AOI22_X1 U1607 ( .A1(reg_mem[501]), .A2(n2896), .B1(n7476), .B2(data_w[5]), 
        .ZN(n2901) );
  INV_X1 U1608 ( .A(n2902), .ZN(n7474) );
  AOI22_X1 U1609 ( .A1(reg_mem[502]), .A2(n2896), .B1(n7476), .B2(data_w[6]), 
        .ZN(n2902) );
  INV_X1 U1610 ( .A(n2903), .ZN(n7475) );
  AOI22_X1 U1611 ( .A1(reg_mem[503]), .A2(n2896), .B1(n7476), .B2(data_w[7]), 
        .ZN(n2903) );
  INV_X1 U1612 ( .A(n2904), .ZN(n8045) );
  AOI22_X1 U1613 ( .A1(reg_mem[504]), .A2(n2905), .B1(n8053), .B2(data_w[0]), 
        .ZN(n2904) );
  INV_X1 U1614 ( .A(n2906), .ZN(n8046) );
  AOI22_X1 U1615 ( .A1(reg_mem[505]), .A2(n2905), .B1(n8053), .B2(data_w[1]), 
        .ZN(n2906) );
  INV_X1 U1616 ( .A(n2907), .ZN(n8047) );
  AOI22_X1 U1617 ( .A1(reg_mem[506]), .A2(n2905), .B1(n8053), .B2(data_w[2]), 
        .ZN(n2907) );
  INV_X1 U1618 ( .A(n2908), .ZN(n8048) );
  AOI22_X1 U1619 ( .A1(reg_mem[507]), .A2(n2905), .B1(n8053), .B2(data_w[3]), 
        .ZN(n2908) );
  INV_X1 U1620 ( .A(n2909), .ZN(n8049) );
  AOI22_X1 U1621 ( .A1(reg_mem[508]), .A2(n2905), .B1(n8053), .B2(data_w[4]), 
        .ZN(n2909) );
  INV_X1 U1622 ( .A(n2910), .ZN(n8050) );
  AOI22_X1 U1623 ( .A1(reg_mem[509]), .A2(n2905), .B1(n8053), .B2(data_w[5]), 
        .ZN(n2910) );
  INV_X1 U1624 ( .A(n2911), .ZN(n8051) );
  AOI22_X1 U1625 ( .A1(reg_mem[510]), .A2(n2905), .B1(n8053), .B2(data_w[6]), 
        .ZN(n2911) );
  INV_X1 U1626 ( .A(n2912), .ZN(n8052) );
  AOI22_X1 U1627 ( .A1(reg_mem[511]), .A2(n2905), .B1(n8053), .B2(data_w[7]), 
        .ZN(n2912) );
  INV_X1 U1628 ( .A(n2914), .ZN(n7315) );
  AOI22_X1 U1629 ( .A1(reg_mem[512]), .A2(n2915), .B1(n7323), .B2(data_w[0]), 
        .ZN(n2914) );
  INV_X1 U1630 ( .A(n2916), .ZN(n7316) );
  AOI22_X1 U1631 ( .A1(reg_mem[513]), .A2(n2915), .B1(n7323), .B2(data_w[1]), 
        .ZN(n2916) );
  INV_X1 U1632 ( .A(n2917), .ZN(n7317) );
  AOI22_X1 U1633 ( .A1(reg_mem[514]), .A2(n2915), .B1(n7323), .B2(data_w[2]), 
        .ZN(n2917) );
  INV_X1 U1634 ( .A(n2918), .ZN(n7318) );
  AOI22_X1 U1635 ( .A1(reg_mem[515]), .A2(n2915), .B1(n7323), .B2(data_w[3]), 
        .ZN(n2918) );
  INV_X1 U1636 ( .A(n2919), .ZN(n7319) );
  AOI22_X1 U1637 ( .A1(reg_mem[516]), .A2(n2915), .B1(n7323), .B2(data_w[4]), 
        .ZN(n2919) );
  INV_X1 U1638 ( .A(n2920), .ZN(n7320) );
  AOI22_X1 U1639 ( .A1(reg_mem[517]), .A2(n2915), .B1(n7323), .B2(data_w[5]), 
        .ZN(n2920) );
  INV_X1 U1640 ( .A(n2921), .ZN(n7321) );
  AOI22_X1 U1641 ( .A1(reg_mem[518]), .A2(n2915), .B1(n7323), .B2(data_w[6]), 
        .ZN(n2921) );
  INV_X1 U1642 ( .A(n2922), .ZN(n7322) );
  AOI22_X1 U1643 ( .A1(reg_mem[519]), .A2(n2915), .B1(n7323), .B2(data_w[7]), 
        .ZN(n2922) );
  INV_X1 U1644 ( .A(n2924), .ZN(n9044) );
  AOI22_X1 U1645 ( .A1(reg_mem[520]), .A2(n2925), .B1(n9052), .B2(data_w[0]), 
        .ZN(n2924) );
  INV_X1 U1646 ( .A(n2926), .ZN(n9045) );
  AOI22_X1 U1647 ( .A1(reg_mem[521]), .A2(n2925), .B1(n9052), .B2(data_w[1]), 
        .ZN(n2926) );
  INV_X1 U1648 ( .A(n2927), .ZN(n9046) );
  AOI22_X1 U1649 ( .A1(reg_mem[522]), .A2(n2925), .B1(n9052), .B2(data_w[2]), 
        .ZN(n2927) );
  INV_X1 U1650 ( .A(n2928), .ZN(n9047) );
  AOI22_X1 U1651 ( .A1(reg_mem[523]), .A2(n2925), .B1(n9052), .B2(data_w[3]), 
        .ZN(n2928) );
  INV_X1 U1652 ( .A(n2929), .ZN(n9048) );
  AOI22_X1 U1653 ( .A1(reg_mem[524]), .A2(n2925), .B1(n9052), .B2(data_w[4]), 
        .ZN(n2929) );
  INV_X1 U1654 ( .A(n2930), .ZN(n9049) );
  AOI22_X1 U1655 ( .A1(reg_mem[525]), .A2(n2925), .B1(n9052), .B2(data_w[5]), 
        .ZN(n2930) );
  INV_X1 U1656 ( .A(n2931), .ZN(n9050) );
  AOI22_X1 U1657 ( .A1(reg_mem[526]), .A2(n2925), .B1(n9052), .B2(data_w[6]), 
        .ZN(n2931) );
  INV_X1 U1658 ( .A(n2932), .ZN(n9051) );
  AOI22_X1 U1659 ( .A1(reg_mem[527]), .A2(n2925), .B1(n9052), .B2(data_w[7]), 
        .ZN(n2932) );
  INV_X1 U1660 ( .A(n2933), .ZN(n7891) );
  AOI22_X1 U1661 ( .A1(reg_mem[528]), .A2(n2934), .B1(n7899), .B2(data_w[0]), 
        .ZN(n2933) );
  INV_X1 U1662 ( .A(n2935), .ZN(n7892) );
  AOI22_X1 U1663 ( .A1(reg_mem[529]), .A2(n2934), .B1(n7899), .B2(data_w[1]), 
        .ZN(n2935) );
  INV_X1 U1664 ( .A(n2936), .ZN(n7893) );
  AOI22_X1 U1665 ( .A1(reg_mem[530]), .A2(n2934), .B1(n7899), .B2(data_w[2]), 
        .ZN(n2936) );
  INV_X1 U1666 ( .A(n2937), .ZN(n7894) );
  AOI22_X1 U1667 ( .A1(reg_mem[531]), .A2(n2934), .B1(n7899), .B2(data_w[3]), 
        .ZN(n2937) );
  INV_X1 U1668 ( .A(n2938), .ZN(n7895) );
  AOI22_X1 U1669 ( .A1(reg_mem[532]), .A2(n2934), .B1(n7899), .B2(data_w[4]), 
        .ZN(n2938) );
  INV_X1 U1670 ( .A(n2939), .ZN(n7896) );
  AOI22_X1 U1671 ( .A1(reg_mem[533]), .A2(n2934), .B1(n7899), .B2(data_w[5]), 
        .ZN(n2939) );
  INV_X1 U1672 ( .A(n2940), .ZN(n7897) );
  AOI22_X1 U1673 ( .A1(reg_mem[534]), .A2(n2934), .B1(n7899), .B2(data_w[6]), 
        .ZN(n2940) );
  INV_X1 U1674 ( .A(n2941), .ZN(n7898) );
  AOI22_X1 U1675 ( .A1(reg_mem[535]), .A2(n2934), .B1(n7899), .B2(data_w[7]), 
        .ZN(n2941) );
  INV_X1 U1676 ( .A(n2942), .ZN(n8468) );
  AOI22_X1 U1677 ( .A1(reg_mem[536]), .A2(n2943), .B1(n8476), .B2(data_w[0]), 
        .ZN(n2942) );
  INV_X1 U1678 ( .A(n2944), .ZN(n8469) );
  AOI22_X1 U1679 ( .A1(reg_mem[537]), .A2(n2943), .B1(n8476), .B2(data_w[1]), 
        .ZN(n2944) );
  INV_X1 U1680 ( .A(n2945), .ZN(n8470) );
  AOI22_X1 U1681 ( .A1(reg_mem[538]), .A2(n2943), .B1(n8476), .B2(data_w[2]), 
        .ZN(n2945) );
  INV_X1 U1682 ( .A(n2946), .ZN(n8471) );
  AOI22_X1 U1683 ( .A1(reg_mem[539]), .A2(n2943), .B1(n8476), .B2(data_w[3]), 
        .ZN(n2946) );
  INV_X1 U1684 ( .A(n2947), .ZN(n8472) );
  AOI22_X1 U1685 ( .A1(reg_mem[540]), .A2(n2943), .B1(n8476), .B2(data_w[4]), 
        .ZN(n2947) );
  INV_X1 U1686 ( .A(n2948), .ZN(n8473) );
  AOI22_X1 U1687 ( .A1(reg_mem[541]), .A2(n2943), .B1(n8476), .B2(data_w[5]), 
        .ZN(n2948) );
  INV_X1 U1688 ( .A(n2949), .ZN(n8474) );
  AOI22_X1 U1689 ( .A1(reg_mem[542]), .A2(n2943), .B1(n8476), .B2(data_w[6]), 
        .ZN(n2949) );
  INV_X1 U1690 ( .A(n2950), .ZN(n8475) );
  AOI22_X1 U1691 ( .A1(reg_mem[543]), .A2(n2943), .B1(n8476), .B2(data_w[7]), 
        .ZN(n2950) );
  INV_X1 U1692 ( .A(n2951), .ZN(n7171) );
  AOI22_X1 U1693 ( .A1(reg_mem[544]), .A2(n2952), .B1(n7179), .B2(data_w[0]), 
        .ZN(n2951) );
  INV_X1 U1694 ( .A(n2953), .ZN(n7172) );
  AOI22_X1 U1695 ( .A1(reg_mem[545]), .A2(n2952), .B1(n7179), .B2(data_w[1]), 
        .ZN(n2953) );
  INV_X1 U1696 ( .A(n2954), .ZN(n7173) );
  AOI22_X1 U1697 ( .A1(reg_mem[546]), .A2(n2952), .B1(n7179), .B2(data_w[2]), 
        .ZN(n2954) );
  INV_X1 U1698 ( .A(n2955), .ZN(n7174) );
  AOI22_X1 U1699 ( .A1(reg_mem[547]), .A2(n2952), .B1(n7179), .B2(data_w[3]), 
        .ZN(n2955) );
  INV_X1 U1700 ( .A(n2956), .ZN(n7175) );
  AOI22_X1 U1701 ( .A1(reg_mem[548]), .A2(n2952), .B1(n7179), .B2(data_w[4]), 
        .ZN(n2956) );
  INV_X1 U1702 ( .A(n2957), .ZN(n7176) );
  AOI22_X1 U1703 ( .A1(reg_mem[549]), .A2(n2952), .B1(n7179), .B2(data_w[5]), 
        .ZN(n2957) );
  INV_X1 U1704 ( .A(n2958), .ZN(n7177) );
  AOI22_X1 U1705 ( .A1(reg_mem[550]), .A2(n2952), .B1(n7179), .B2(data_w[6]), 
        .ZN(n2958) );
  INV_X1 U1706 ( .A(n2959), .ZN(n7178) );
  AOI22_X1 U1707 ( .A1(reg_mem[551]), .A2(n2952), .B1(n7179), .B2(data_w[7]), 
        .ZN(n2959) );
  INV_X1 U1708 ( .A(n2960), .ZN(n8900) );
  AOI22_X1 U1709 ( .A1(reg_mem[552]), .A2(n2961), .B1(n8908), .B2(data_w[0]), 
        .ZN(n2960) );
  INV_X1 U1710 ( .A(n2962), .ZN(n8901) );
  AOI22_X1 U1711 ( .A1(reg_mem[553]), .A2(n2961), .B1(n8908), .B2(data_w[1]), 
        .ZN(n2962) );
  INV_X1 U1712 ( .A(n2963), .ZN(n8902) );
  AOI22_X1 U1713 ( .A1(reg_mem[554]), .A2(n2961), .B1(n8908), .B2(data_w[2]), 
        .ZN(n2963) );
  INV_X1 U1714 ( .A(n2964), .ZN(n8903) );
  AOI22_X1 U1715 ( .A1(reg_mem[555]), .A2(n2961), .B1(n8908), .B2(data_w[3]), 
        .ZN(n2964) );
  INV_X1 U1716 ( .A(n2965), .ZN(n8904) );
  AOI22_X1 U1717 ( .A1(reg_mem[556]), .A2(n2961), .B1(n8908), .B2(data_w[4]), 
        .ZN(n2965) );
  INV_X1 U1718 ( .A(n2966), .ZN(n8905) );
  AOI22_X1 U1719 ( .A1(reg_mem[557]), .A2(n2961), .B1(n8908), .B2(data_w[5]), 
        .ZN(n2966) );
  INV_X1 U1720 ( .A(n2967), .ZN(n8906) );
  AOI22_X1 U1721 ( .A1(reg_mem[558]), .A2(n2961), .B1(n8908), .B2(data_w[6]), 
        .ZN(n2967) );
  INV_X1 U1722 ( .A(n2968), .ZN(n8907) );
  AOI22_X1 U1723 ( .A1(reg_mem[559]), .A2(n2961), .B1(n8908), .B2(data_w[7]), 
        .ZN(n2968) );
  INV_X1 U1724 ( .A(n2969), .ZN(n7747) );
  AOI22_X1 U1725 ( .A1(reg_mem[560]), .A2(n2970), .B1(n7755), .B2(data_w[0]), 
        .ZN(n2969) );
  INV_X1 U1726 ( .A(n2971), .ZN(n7748) );
  AOI22_X1 U1727 ( .A1(reg_mem[561]), .A2(n2970), .B1(n7755), .B2(data_w[1]), 
        .ZN(n2971) );
  INV_X1 U1728 ( .A(n2972), .ZN(n7749) );
  AOI22_X1 U1729 ( .A1(reg_mem[562]), .A2(n2970), .B1(n7755), .B2(data_w[2]), 
        .ZN(n2972) );
  INV_X1 U1730 ( .A(n2973), .ZN(n7750) );
  AOI22_X1 U1731 ( .A1(reg_mem[563]), .A2(n2970), .B1(n7755), .B2(data_w[3]), 
        .ZN(n2973) );
  INV_X1 U1732 ( .A(n2974), .ZN(n7751) );
  AOI22_X1 U1733 ( .A1(reg_mem[564]), .A2(n2970), .B1(n7755), .B2(data_w[4]), 
        .ZN(n2974) );
  INV_X1 U1734 ( .A(n2975), .ZN(n7752) );
  AOI22_X1 U1735 ( .A1(reg_mem[565]), .A2(n2970), .B1(n7755), .B2(data_w[5]), 
        .ZN(n2975) );
  INV_X1 U1736 ( .A(n2976), .ZN(n7753) );
  AOI22_X1 U1737 ( .A1(reg_mem[566]), .A2(n2970), .B1(n7755), .B2(data_w[6]), 
        .ZN(n2976) );
  INV_X1 U1738 ( .A(n2977), .ZN(n7754) );
  AOI22_X1 U1739 ( .A1(reg_mem[567]), .A2(n2970), .B1(n7755), .B2(data_w[7]), 
        .ZN(n2977) );
  INV_X1 U1740 ( .A(n2978), .ZN(n8324) );
  AOI22_X1 U1741 ( .A1(reg_mem[568]), .A2(n2979), .B1(n8332), .B2(data_w[0]), 
        .ZN(n2978) );
  INV_X1 U1742 ( .A(n2980), .ZN(n8325) );
  AOI22_X1 U1743 ( .A1(reg_mem[569]), .A2(n2979), .B1(n8332), .B2(data_w[1]), 
        .ZN(n2980) );
  INV_X1 U1744 ( .A(n2981), .ZN(n8326) );
  AOI22_X1 U1745 ( .A1(reg_mem[570]), .A2(n2979), .B1(n8332), .B2(data_w[2]), 
        .ZN(n2981) );
  INV_X1 U1746 ( .A(n2982), .ZN(n8327) );
  AOI22_X1 U1747 ( .A1(reg_mem[571]), .A2(n2979), .B1(n8332), .B2(data_w[3]), 
        .ZN(n2982) );
  INV_X1 U1748 ( .A(n2983), .ZN(n8328) );
  AOI22_X1 U1749 ( .A1(reg_mem[572]), .A2(n2979), .B1(n8332), .B2(data_w[4]), 
        .ZN(n2983) );
  INV_X1 U1750 ( .A(n2984), .ZN(n8329) );
  AOI22_X1 U1751 ( .A1(reg_mem[573]), .A2(n2979), .B1(n8332), .B2(data_w[5]), 
        .ZN(n2984) );
  INV_X1 U1752 ( .A(n2985), .ZN(n8330) );
  AOI22_X1 U1753 ( .A1(reg_mem[574]), .A2(n2979), .B1(n8332), .B2(data_w[6]), 
        .ZN(n2985) );
  INV_X1 U1754 ( .A(n2986), .ZN(n8331) );
  AOI22_X1 U1755 ( .A1(reg_mem[575]), .A2(n2979), .B1(n8332), .B2(data_w[7]), 
        .ZN(n2986) );
  INV_X1 U1756 ( .A(n2987), .ZN(n7027) );
  AOI22_X1 U1757 ( .A1(reg_mem[576]), .A2(n2988), .B1(n7035), .B2(data_w[0]), 
        .ZN(n2987) );
  INV_X1 U1758 ( .A(n2989), .ZN(n7028) );
  AOI22_X1 U1759 ( .A1(reg_mem[577]), .A2(n2988), .B1(n7035), .B2(data_w[1]), 
        .ZN(n2989) );
  INV_X1 U1760 ( .A(n2990), .ZN(n7029) );
  AOI22_X1 U1761 ( .A1(reg_mem[578]), .A2(n2988), .B1(n7035), .B2(data_w[2]), 
        .ZN(n2990) );
  INV_X1 U1762 ( .A(n2991), .ZN(n7030) );
  AOI22_X1 U1763 ( .A1(reg_mem[579]), .A2(n2988), .B1(n7035), .B2(data_w[3]), 
        .ZN(n2991) );
  INV_X1 U1764 ( .A(n2992), .ZN(n7031) );
  AOI22_X1 U1765 ( .A1(reg_mem[580]), .A2(n2988), .B1(n7035), .B2(data_w[4]), 
        .ZN(n2992) );
  INV_X1 U1766 ( .A(n2993), .ZN(n7032) );
  AOI22_X1 U1767 ( .A1(reg_mem[581]), .A2(n2988), .B1(n7035), .B2(data_w[5]), 
        .ZN(n2993) );
  INV_X1 U1768 ( .A(n2994), .ZN(n7033) );
  AOI22_X1 U1769 ( .A1(reg_mem[582]), .A2(n2988), .B1(n7035), .B2(data_w[6]), 
        .ZN(n2994) );
  INV_X1 U1770 ( .A(n2995), .ZN(n7034) );
  AOI22_X1 U1771 ( .A1(reg_mem[583]), .A2(n2988), .B1(n7035), .B2(data_w[7]), 
        .ZN(n2995) );
  INV_X1 U1772 ( .A(n2996), .ZN(n8756) );
  AOI22_X1 U1773 ( .A1(reg_mem[584]), .A2(n2997), .B1(n8764), .B2(data_w[0]), 
        .ZN(n2996) );
  INV_X1 U1774 ( .A(n2998), .ZN(n8757) );
  AOI22_X1 U1775 ( .A1(reg_mem[585]), .A2(n2997), .B1(n8764), .B2(data_w[1]), 
        .ZN(n2998) );
  INV_X1 U1776 ( .A(n2999), .ZN(n8758) );
  AOI22_X1 U1777 ( .A1(reg_mem[586]), .A2(n2997), .B1(n8764), .B2(data_w[2]), 
        .ZN(n2999) );
  INV_X1 U1778 ( .A(n3000), .ZN(n8759) );
  AOI22_X1 U1779 ( .A1(reg_mem[587]), .A2(n2997), .B1(n8764), .B2(data_w[3]), 
        .ZN(n3000) );
  INV_X1 U1780 ( .A(n3001), .ZN(n8760) );
  AOI22_X1 U1781 ( .A1(reg_mem[588]), .A2(n2997), .B1(n8764), .B2(data_w[4]), 
        .ZN(n3001) );
  INV_X1 U1782 ( .A(n3002), .ZN(n8761) );
  AOI22_X1 U1783 ( .A1(reg_mem[589]), .A2(n2997), .B1(n8764), .B2(data_w[5]), 
        .ZN(n3002) );
  INV_X1 U1784 ( .A(n3003), .ZN(n8762) );
  AOI22_X1 U1785 ( .A1(reg_mem[590]), .A2(n2997), .B1(n8764), .B2(data_w[6]), 
        .ZN(n3003) );
  INV_X1 U1786 ( .A(n3004), .ZN(n8763) );
  AOI22_X1 U1787 ( .A1(reg_mem[591]), .A2(n2997), .B1(n8764), .B2(data_w[7]), 
        .ZN(n3004) );
  INV_X1 U1788 ( .A(n3005), .ZN(n7603) );
  AOI22_X1 U1789 ( .A1(reg_mem[592]), .A2(n3006), .B1(n7611), .B2(data_w[0]), 
        .ZN(n3005) );
  INV_X1 U1790 ( .A(n3007), .ZN(n7604) );
  AOI22_X1 U1791 ( .A1(reg_mem[593]), .A2(n3006), .B1(n7611), .B2(data_w[1]), 
        .ZN(n3007) );
  INV_X1 U1792 ( .A(n3008), .ZN(n7605) );
  AOI22_X1 U1793 ( .A1(reg_mem[594]), .A2(n3006), .B1(n7611), .B2(data_w[2]), 
        .ZN(n3008) );
  INV_X1 U1794 ( .A(n3009), .ZN(n7606) );
  AOI22_X1 U1795 ( .A1(reg_mem[595]), .A2(n3006), .B1(n7611), .B2(data_w[3]), 
        .ZN(n3009) );
  INV_X1 U1796 ( .A(n3010), .ZN(n7607) );
  AOI22_X1 U1797 ( .A1(reg_mem[596]), .A2(n3006), .B1(n7611), .B2(data_w[4]), 
        .ZN(n3010) );
  INV_X1 U1798 ( .A(n3011), .ZN(n7608) );
  AOI22_X1 U1799 ( .A1(reg_mem[597]), .A2(n3006), .B1(n7611), .B2(data_w[5]), 
        .ZN(n3011) );
  INV_X1 U1800 ( .A(n3012), .ZN(n7609) );
  AOI22_X1 U1801 ( .A1(reg_mem[598]), .A2(n3006), .B1(n7611), .B2(data_w[6]), 
        .ZN(n3012) );
  INV_X1 U1802 ( .A(n3013), .ZN(n7610) );
  AOI22_X1 U1803 ( .A1(reg_mem[599]), .A2(n3006), .B1(n7611), .B2(data_w[7]), 
        .ZN(n3013) );
  INV_X1 U1804 ( .A(n3014), .ZN(n8180) );
  AOI22_X1 U1805 ( .A1(reg_mem[600]), .A2(n3015), .B1(n8188), .B2(data_w[0]), 
        .ZN(n3014) );
  INV_X1 U1806 ( .A(n3016), .ZN(n8181) );
  AOI22_X1 U1807 ( .A1(reg_mem[601]), .A2(n3015), .B1(n8188), .B2(data_w[1]), 
        .ZN(n3016) );
  INV_X1 U1808 ( .A(n3017), .ZN(n8182) );
  AOI22_X1 U1809 ( .A1(reg_mem[602]), .A2(n3015), .B1(n8188), .B2(data_w[2]), 
        .ZN(n3017) );
  INV_X1 U1810 ( .A(n3018), .ZN(n8183) );
  AOI22_X1 U1811 ( .A1(reg_mem[603]), .A2(n3015), .B1(n8188), .B2(data_w[3]), 
        .ZN(n3018) );
  INV_X1 U1812 ( .A(n3019), .ZN(n8184) );
  AOI22_X1 U1813 ( .A1(reg_mem[604]), .A2(n3015), .B1(n8188), .B2(data_w[4]), 
        .ZN(n3019) );
  INV_X1 U1814 ( .A(n3020), .ZN(n8185) );
  AOI22_X1 U1815 ( .A1(reg_mem[605]), .A2(n3015), .B1(n8188), .B2(data_w[5]), 
        .ZN(n3020) );
  INV_X1 U1816 ( .A(n3021), .ZN(n8186) );
  AOI22_X1 U1817 ( .A1(reg_mem[606]), .A2(n3015), .B1(n8188), .B2(data_w[6]), 
        .ZN(n3021) );
  INV_X1 U1818 ( .A(n3022), .ZN(n8187) );
  AOI22_X1 U1819 ( .A1(reg_mem[607]), .A2(n3015), .B1(n8188), .B2(data_w[7]), 
        .ZN(n3022) );
  INV_X1 U1820 ( .A(n3023), .ZN(n6883) );
  AOI22_X1 U1821 ( .A1(reg_mem[608]), .A2(n3024), .B1(n6891), .B2(data_w[0]), 
        .ZN(n3023) );
  INV_X1 U1822 ( .A(n3025), .ZN(n6884) );
  AOI22_X1 U1823 ( .A1(reg_mem[609]), .A2(n3024), .B1(n6891), .B2(data_w[1]), 
        .ZN(n3025) );
  INV_X1 U1824 ( .A(n3026), .ZN(n6885) );
  AOI22_X1 U1825 ( .A1(reg_mem[610]), .A2(n3024), .B1(n6891), .B2(data_w[2]), 
        .ZN(n3026) );
  INV_X1 U1826 ( .A(n3027), .ZN(n6886) );
  AOI22_X1 U1827 ( .A1(reg_mem[611]), .A2(n3024), .B1(n6891), .B2(data_w[3]), 
        .ZN(n3027) );
  INV_X1 U1828 ( .A(n3028), .ZN(n6887) );
  AOI22_X1 U1829 ( .A1(reg_mem[612]), .A2(n3024), .B1(n6891), .B2(data_w[4]), 
        .ZN(n3028) );
  INV_X1 U1830 ( .A(n3029), .ZN(n6888) );
  AOI22_X1 U1831 ( .A1(reg_mem[613]), .A2(n3024), .B1(n6891), .B2(data_w[5]), 
        .ZN(n3029) );
  INV_X1 U1832 ( .A(n3030), .ZN(n6889) );
  AOI22_X1 U1833 ( .A1(reg_mem[614]), .A2(n3024), .B1(n6891), .B2(data_w[6]), 
        .ZN(n3030) );
  INV_X1 U1834 ( .A(n3031), .ZN(n6890) );
  AOI22_X1 U1835 ( .A1(reg_mem[615]), .A2(n3024), .B1(n6891), .B2(data_w[7]), 
        .ZN(n3031) );
  INV_X1 U1836 ( .A(n3032), .ZN(n8612) );
  AOI22_X1 U1837 ( .A1(reg_mem[616]), .A2(n3033), .B1(n8620), .B2(data_w[0]), 
        .ZN(n3032) );
  INV_X1 U1838 ( .A(n3034), .ZN(n8613) );
  AOI22_X1 U1839 ( .A1(reg_mem[617]), .A2(n3033), .B1(n8620), .B2(data_w[1]), 
        .ZN(n3034) );
  INV_X1 U1840 ( .A(n3035), .ZN(n8614) );
  AOI22_X1 U1841 ( .A1(reg_mem[618]), .A2(n3033), .B1(n8620), .B2(data_w[2]), 
        .ZN(n3035) );
  INV_X1 U1842 ( .A(n3036), .ZN(n8615) );
  AOI22_X1 U1843 ( .A1(reg_mem[619]), .A2(n3033), .B1(n8620), .B2(data_w[3]), 
        .ZN(n3036) );
  INV_X1 U1844 ( .A(n3037), .ZN(n8616) );
  AOI22_X1 U1845 ( .A1(reg_mem[620]), .A2(n3033), .B1(n8620), .B2(data_w[4]), 
        .ZN(n3037) );
  INV_X1 U1846 ( .A(n3038), .ZN(n8617) );
  AOI22_X1 U1847 ( .A1(reg_mem[621]), .A2(n3033), .B1(n8620), .B2(data_w[5]), 
        .ZN(n3038) );
  INV_X1 U1848 ( .A(n3039), .ZN(n8618) );
  AOI22_X1 U1849 ( .A1(reg_mem[622]), .A2(n3033), .B1(n8620), .B2(data_w[6]), 
        .ZN(n3039) );
  INV_X1 U1850 ( .A(n3040), .ZN(n8619) );
  AOI22_X1 U1851 ( .A1(reg_mem[623]), .A2(n3033), .B1(n8620), .B2(data_w[7]), 
        .ZN(n3040) );
  INV_X1 U1852 ( .A(n3041), .ZN(n7459) );
  AOI22_X1 U1853 ( .A1(reg_mem[624]), .A2(n3042), .B1(n7467), .B2(data_w[0]), 
        .ZN(n3041) );
  INV_X1 U1854 ( .A(n3043), .ZN(n7460) );
  AOI22_X1 U1855 ( .A1(reg_mem[625]), .A2(n3042), .B1(n7467), .B2(data_w[1]), 
        .ZN(n3043) );
  INV_X1 U1856 ( .A(n3044), .ZN(n7461) );
  AOI22_X1 U1857 ( .A1(reg_mem[626]), .A2(n3042), .B1(n7467), .B2(data_w[2]), 
        .ZN(n3044) );
  INV_X1 U1858 ( .A(n3045), .ZN(n7462) );
  AOI22_X1 U1859 ( .A1(reg_mem[627]), .A2(n3042), .B1(n7467), .B2(data_w[3]), 
        .ZN(n3045) );
  INV_X1 U1860 ( .A(n3046), .ZN(n7463) );
  AOI22_X1 U1861 ( .A1(reg_mem[628]), .A2(n3042), .B1(n7467), .B2(data_w[4]), 
        .ZN(n3046) );
  INV_X1 U1862 ( .A(n3047), .ZN(n7464) );
  AOI22_X1 U1863 ( .A1(reg_mem[629]), .A2(n3042), .B1(n7467), .B2(data_w[5]), 
        .ZN(n3047) );
  INV_X1 U1864 ( .A(n3048), .ZN(n7465) );
  AOI22_X1 U1865 ( .A1(reg_mem[630]), .A2(n3042), .B1(n7467), .B2(data_w[6]), 
        .ZN(n3048) );
  INV_X1 U1866 ( .A(n3049), .ZN(n7466) );
  AOI22_X1 U1867 ( .A1(reg_mem[631]), .A2(n3042), .B1(n7467), .B2(data_w[7]), 
        .ZN(n3049) );
  INV_X1 U1868 ( .A(n3050), .ZN(n8036) );
  AOI22_X1 U1869 ( .A1(reg_mem[632]), .A2(n3051), .B1(n8044), .B2(data_w[0]), 
        .ZN(n3050) );
  INV_X1 U1870 ( .A(n3052), .ZN(n8037) );
  AOI22_X1 U1871 ( .A1(reg_mem[633]), .A2(n3051), .B1(n8044), .B2(data_w[1]), 
        .ZN(n3052) );
  INV_X1 U1872 ( .A(n3053), .ZN(n8038) );
  AOI22_X1 U1873 ( .A1(reg_mem[634]), .A2(n3051), .B1(n8044), .B2(data_w[2]), 
        .ZN(n3053) );
  INV_X1 U1874 ( .A(n3054), .ZN(n8039) );
  AOI22_X1 U1875 ( .A1(reg_mem[635]), .A2(n3051), .B1(n8044), .B2(data_w[3]), 
        .ZN(n3054) );
  INV_X1 U1876 ( .A(n3055), .ZN(n8040) );
  AOI22_X1 U1877 ( .A1(reg_mem[636]), .A2(n3051), .B1(n8044), .B2(data_w[4]), 
        .ZN(n3055) );
  INV_X1 U1878 ( .A(n3056), .ZN(n8041) );
  AOI22_X1 U1879 ( .A1(reg_mem[637]), .A2(n3051), .B1(n8044), .B2(data_w[5]), 
        .ZN(n3056) );
  INV_X1 U1880 ( .A(n3057), .ZN(n8042) );
  AOI22_X1 U1881 ( .A1(reg_mem[638]), .A2(n3051), .B1(n8044), .B2(data_w[6]), 
        .ZN(n3057) );
  INV_X1 U1882 ( .A(n3058), .ZN(n8043) );
  AOI22_X1 U1883 ( .A1(reg_mem[639]), .A2(n3051), .B1(n8044), .B2(data_w[7]), 
        .ZN(n3058) );
  INV_X1 U1884 ( .A(n3060), .ZN(n7306) );
  AOI22_X1 U1885 ( .A1(reg_mem[640]), .A2(n3061), .B1(n7314), .B2(data_w[0]), 
        .ZN(n3060) );
  INV_X1 U1886 ( .A(n3062), .ZN(n7307) );
  AOI22_X1 U1887 ( .A1(reg_mem[641]), .A2(n3061), .B1(n7314), .B2(data_w[1]), 
        .ZN(n3062) );
  INV_X1 U1888 ( .A(n3063), .ZN(n7308) );
  AOI22_X1 U1889 ( .A1(reg_mem[642]), .A2(n3061), .B1(n7314), .B2(data_w[2]), 
        .ZN(n3063) );
  INV_X1 U1890 ( .A(n3064), .ZN(n7309) );
  AOI22_X1 U1891 ( .A1(reg_mem[643]), .A2(n3061), .B1(n7314), .B2(data_w[3]), 
        .ZN(n3064) );
  INV_X1 U1892 ( .A(n3065), .ZN(n7310) );
  AOI22_X1 U1893 ( .A1(reg_mem[644]), .A2(n3061), .B1(n7314), .B2(data_w[4]), 
        .ZN(n3065) );
  INV_X1 U1894 ( .A(n3066), .ZN(n7311) );
  AOI22_X1 U1895 ( .A1(reg_mem[645]), .A2(n3061), .B1(n7314), .B2(data_w[5]), 
        .ZN(n3066) );
  INV_X1 U1896 ( .A(n3067), .ZN(n7312) );
  AOI22_X1 U1897 ( .A1(reg_mem[646]), .A2(n3061), .B1(n7314), .B2(data_w[6]), 
        .ZN(n3067) );
  INV_X1 U1898 ( .A(n3068), .ZN(n7313) );
  AOI22_X1 U1899 ( .A1(reg_mem[647]), .A2(n3061), .B1(n7314), .B2(data_w[7]), 
        .ZN(n3068) );
  INV_X1 U1900 ( .A(n3070), .ZN(n9035) );
  AOI22_X1 U1901 ( .A1(reg_mem[648]), .A2(n3071), .B1(n9043), .B2(data_w[0]), 
        .ZN(n3070) );
  INV_X1 U1902 ( .A(n3072), .ZN(n9036) );
  AOI22_X1 U1903 ( .A1(reg_mem[649]), .A2(n3071), .B1(n9043), .B2(data_w[1]), 
        .ZN(n3072) );
  INV_X1 U1904 ( .A(n3073), .ZN(n9037) );
  AOI22_X1 U1905 ( .A1(reg_mem[650]), .A2(n3071), .B1(n9043), .B2(data_w[2]), 
        .ZN(n3073) );
  INV_X1 U1906 ( .A(n3074), .ZN(n9038) );
  AOI22_X1 U1907 ( .A1(reg_mem[651]), .A2(n3071), .B1(n9043), .B2(data_w[3]), 
        .ZN(n3074) );
  INV_X1 U1908 ( .A(n3075), .ZN(n9039) );
  AOI22_X1 U1909 ( .A1(reg_mem[652]), .A2(n3071), .B1(n9043), .B2(data_w[4]), 
        .ZN(n3075) );
  INV_X1 U1910 ( .A(n3076), .ZN(n9040) );
  AOI22_X1 U1911 ( .A1(reg_mem[653]), .A2(n3071), .B1(n9043), .B2(data_w[5]), 
        .ZN(n3076) );
  INV_X1 U1912 ( .A(n3077), .ZN(n9041) );
  AOI22_X1 U1913 ( .A1(reg_mem[654]), .A2(n3071), .B1(n9043), .B2(data_w[6]), 
        .ZN(n3077) );
  INV_X1 U1914 ( .A(n3078), .ZN(n9042) );
  AOI22_X1 U1915 ( .A1(reg_mem[655]), .A2(n3071), .B1(n9043), .B2(data_w[7]), 
        .ZN(n3078) );
  INV_X1 U1916 ( .A(n3079), .ZN(n7882) );
  AOI22_X1 U1917 ( .A1(reg_mem[656]), .A2(n3080), .B1(n7890), .B2(data_w[0]), 
        .ZN(n3079) );
  INV_X1 U1918 ( .A(n3081), .ZN(n7883) );
  AOI22_X1 U1919 ( .A1(reg_mem[657]), .A2(n3080), .B1(n7890), .B2(data_w[1]), 
        .ZN(n3081) );
  INV_X1 U1920 ( .A(n3082), .ZN(n7884) );
  AOI22_X1 U1921 ( .A1(reg_mem[658]), .A2(n3080), .B1(n7890), .B2(data_w[2]), 
        .ZN(n3082) );
  INV_X1 U1922 ( .A(n3083), .ZN(n7885) );
  AOI22_X1 U1923 ( .A1(reg_mem[659]), .A2(n3080), .B1(n7890), .B2(data_w[3]), 
        .ZN(n3083) );
  INV_X1 U1924 ( .A(n3084), .ZN(n7886) );
  AOI22_X1 U1925 ( .A1(reg_mem[660]), .A2(n3080), .B1(n7890), .B2(data_w[4]), 
        .ZN(n3084) );
  INV_X1 U1926 ( .A(n3085), .ZN(n7887) );
  AOI22_X1 U1927 ( .A1(reg_mem[661]), .A2(n3080), .B1(n7890), .B2(data_w[5]), 
        .ZN(n3085) );
  INV_X1 U1928 ( .A(n3086), .ZN(n7888) );
  AOI22_X1 U1929 ( .A1(reg_mem[662]), .A2(n3080), .B1(n7890), .B2(data_w[6]), 
        .ZN(n3086) );
  INV_X1 U1930 ( .A(n3087), .ZN(n7889) );
  AOI22_X1 U1931 ( .A1(reg_mem[663]), .A2(n3080), .B1(n7890), .B2(data_w[7]), 
        .ZN(n3087) );
  INV_X1 U1932 ( .A(n3088), .ZN(n8459) );
  AOI22_X1 U1933 ( .A1(reg_mem[664]), .A2(n3089), .B1(n8467), .B2(data_w[0]), 
        .ZN(n3088) );
  INV_X1 U1934 ( .A(n3090), .ZN(n8460) );
  AOI22_X1 U1935 ( .A1(reg_mem[665]), .A2(n3089), .B1(n8467), .B2(data_w[1]), 
        .ZN(n3090) );
  INV_X1 U1936 ( .A(n3091), .ZN(n8461) );
  AOI22_X1 U1937 ( .A1(reg_mem[666]), .A2(n3089), .B1(n8467), .B2(data_w[2]), 
        .ZN(n3091) );
  INV_X1 U1938 ( .A(n3092), .ZN(n8462) );
  AOI22_X1 U1939 ( .A1(reg_mem[667]), .A2(n3089), .B1(n8467), .B2(data_w[3]), 
        .ZN(n3092) );
  INV_X1 U1940 ( .A(n3093), .ZN(n8463) );
  AOI22_X1 U1941 ( .A1(reg_mem[668]), .A2(n3089), .B1(n8467), .B2(data_w[4]), 
        .ZN(n3093) );
  INV_X1 U1942 ( .A(n3094), .ZN(n8464) );
  AOI22_X1 U1943 ( .A1(reg_mem[669]), .A2(n3089), .B1(n8467), .B2(data_w[5]), 
        .ZN(n3094) );
  INV_X1 U1944 ( .A(n3095), .ZN(n8465) );
  AOI22_X1 U1945 ( .A1(reg_mem[670]), .A2(n3089), .B1(n8467), .B2(data_w[6]), 
        .ZN(n3095) );
  INV_X1 U1946 ( .A(n3096), .ZN(n8466) );
  AOI22_X1 U1947 ( .A1(reg_mem[671]), .A2(n3089), .B1(n8467), .B2(data_w[7]), 
        .ZN(n3096) );
  INV_X1 U1948 ( .A(n3097), .ZN(n7162) );
  AOI22_X1 U1949 ( .A1(reg_mem[672]), .A2(n3098), .B1(n7170), .B2(data_w[0]), 
        .ZN(n3097) );
  INV_X1 U1950 ( .A(n3099), .ZN(n7163) );
  AOI22_X1 U1951 ( .A1(reg_mem[673]), .A2(n3098), .B1(n7170), .B2(data_w[1]), 
        .ZN(n3099) );
  INV_X1 U1952 ( .A(n3100), .ZN(n7164) );
  AOI22_X1 U1953 ( .A1(reg_mem[674]), .A2(n3098), .B1(n7170), .B2(data_w[2]), 
        .ZN(n3100) );
  INV_X1 U1954 ( .A(n3101), .ZN(n7165) );
  AOI22_X1 U1955 ( .A1(reg_mem[675]), .A2(n3098), .B1(n7170), .B2(data_w[3]), 
        .ZN(n3101) );
  INV_X1 U1956 ( .A(n3102), .ZN(n7166) );
  AOI22_X1 U1957 ( .A1(reg_mem[676]), .A2(n3098), .B1(n7170), .B2(data_w[4]), 
        .ZN(n3102) );
  INV_X1 U1958 ( .A(n3103), .ZN(n7167) );
  AOI22_X1 U1959 ( .A1(reg_mem[677]), .A2(n3098), .B1(n7170), .B2(data_w[5]), 
        .ZN(n3103) );
  INV_X1 U1960 ( .A(n3104), .ZN(n7168) );
  AOI22_X1 U1961 ( .A1(reg_mem[678]), .A2(n3098), .B1(n7170), .B2(data_w[6]), 
        .ZN(n3104) );
  INV_X1 U1962 ( .A(n3105), .ZN(n7169) );
  AOI22_X1 U1963 ( .A1(reg_mem[679]), .A2(n3098), .B1(n7170), .B2(data_w[7]), 
        .ZN(n3105) );
  INV_X1 U1964 ( .A(n3106), .ZN(n8891) );
  AOI22_X1 U1965 ( .A1(reg_mem[680]), .A2(n3107), .B1(n8899), .B2(data_w[0]), 
        .ZN(n3106) );
  INV_X1 U1966 ( .A(n3108), .ZN(n8892) );
  AOI22_X1 U1967 ( .A1(reg_mem[681]), .A2(n3107), .B1(n8899), .B2(data_w[1]), 
        .ZN(n3108) );
  INV_X1 U1968 ( .A(n3109), .ZN(n8893) );
  AOI22_X1 U1969 ( .A1(reg_mem[682]), .A2(n3107), .B1(n8899), .B2(data_w[2]), 
        .ZN(n3109) );
  INV_X1 U1970 ( .A(n3110), .ZN(n8894) );
  AOI22_X1 U1971 ( .A1(reg_mem[683]), .A2(n3107), .B1(n8899), .B2(data_w[3]), 
        .ZN(n3110) );
  INV_X1 U1972 ( .A(n3111), .ZN(n8895) );
  AOI22_X1 U1973 ( .A1(reg_mem[684]), .A2(n3107), .B1(n8899), .B2(data_w[4]), 
        .ZN(n3111) );
  INV_X1 U1974 ( .A(n3112), .ZN(n8896) );
  AOI22_X1 U1975 ( .A1(reg_mem[685]), .A2(n3107), .B1(n8899), .B2(data_w[5]), 
        .ZN(n3112) );
  INV_X1 U1976 ( .A(n3113), .ZN(n8897) );
  AOI22_X1 U1977 ( .A1(reg_mem[686]), .A2(n3107), .B1(n8899), .B2(data_w[6]), 
        .ZN(n3113) );
  INV_X1 U1978 ( .A(n3114), .ZN(n8898) );
  AOI22_X1 U1979 ( .A1(reg_mem[687]), .A2(n3107), .B1(n8899), .B2(data_w[7]), 
        .ZN(n3114) );
  INV_X1 U1980 ( .A(n3115), .ZN(n7738) );
  AOI22_X1 U1981 ( .A1(reg_mem[688]), .A2(n3116), .B1(n7746), .B2(data_w[0]), 
        .ZN(n3115) );
  INV_X1 U1982 ( .A(n3117), .ZN(n7739) );
  AOI22_X1 U1983 ( .A1(reg_mem[689]), .A2(n3116), .B1(n7746), .B2(data_w[1]), 
        .ZN(n3117) );
  INV_X1 U1984 ( .A(n3118), .ZN(n7740) );
  AOI22_X1 U1985 ( .A1(reg_mem[690]), .A2(n3116), .B1(n7746), .B2(data_w[2]), 
        .ZN(n3118) );
  INV_X1 U1986 ( .A(n3119), .ZN(n7741) );
  AOI22_X1 U1987 ( .A1(reg_mem[691]), .A2(n3116), .B1(n7746), .B2(data_w[3]), 
        .ZN(n3119) );
  INV_X1 U1988 ( .A(n3120), .ZN(n7742) );
  AOI22_X1 U1989 ( .A1(reg_mem[692]), .A2(n3116), .B1(n7746), .B2(data_w[4]), 
        .ZN(n3120) );
  INV_X1 U1990 ( .A(n3121), .ZN(n7743) );
  AOI22_X1 U1991 ( .A1(reg_mem[693]), .A2(n3116), .B1(n7746), .B2(data_w[5]), 
        .ZN(n3121) );
  INV_X1 U1992 ( .A(n3122), .ZN(n7744) );
  AOI22_X1 U1993 ( .A1(reg_mem[694]), .A2(n3116), .B1(n7746), .B2(data_w[6]), 
        .ZN(n3122) );
  INV_X1 U1994 ( .A(n3123), .ZN(n7745) );
  AOI22_X1 U1995 ( .A1(reg_mem[695]), .A2(n3116), .B1(n7746), .B2(data_w[7]), 
        .ZN(n3123) );
  INV_X1 U1996 ( .A(n3124), .ZN(n8315) );
  AOI22_X1 U1997 ( .A1(reg_mem[696]), .A2(n3125), .B1(n8323), .B2(data_w[0]), 
        .ZN(n3124) );
  INV_X1 U1998 ( .A(n3126), .ZN(n8316) );
  AOI22_X1 U1999 ( .A1(reg_mem[697]), .A2(n3125), .B1(n8323), .B2(data_w[1]), 
        .ZN(n3126) );
  INV_X1 U2000 ( .A(n3127), .ZN(n8317) );
  AOI22_X1 U2001 ( .A1(reg_mem[698]), .A2(n3125), .B1(n8323), .B2(data_w[2]), 
        .ZN(n3127) );
  INV_X1 U2002 ( .A(n3128), .ZN(n8318) );
  AOI22_X1 U2003 ( .A1(reg_mem[699]), .A2(n3125), .B1(n8323), .B2(data_w[3]), 
        .ZN(n3128) );
  INV_X1 U2004 ( .A(n3129), .ZN(n8319) );
  AOI22_X1 U2005 ( .A1(reg_mem[700]), .A2(n3125), .B1(n8323), .B2(data_w[4]), 
        .ZN(n3129) );
  INV_X1 U2006 ( .A(n3130), .ZN(n8320) );
  AOI22_X1 U2007 ( .A1(reg_mem[701]), .A2(n3125), .B1(n8323), .B2(data_w[5]), 
        .ZN(n3130) );
  INV_X1 U2008 ( .A(n3131), .ZN(n8321) );
  AOI22_X1 U2009 ( .A1(reg_mem[702]), .A2(n3125), .B1(n8323), .B2(data_w[6]), 
        .ZN(n3131) );
  INV_X1 U2010 ( .A(n3132), .ZN(n8322) );
  AOI22_X1 U2011 ( .A1(reg_mem[703]), .A2(n3125), .B1(n8323), .B2(data_w[7]), 
        .ZN(n3132) );
  INV_X1 U2012 ( .A(n3133), .ZN(n7018) );
  AOI22_X1 U2013 ( .A1(reg_mem[704]), .A2(n3134), .B1(n7026), .B2(data_w[0]), 
        .ZN(n3133) );
  INV_X1 U2014 ( .A(n3135), .ZN(n7019) );
  AOI22_X1 U2015 ( .A1(reg_mem[705]), .A2(n3134), .B1(n7026), .B2(data_w[1]), 
        .ZN(n3135) );
  INV_X1 U2016 ( .A(n3136), .ZN(n7020) );
  AOI22_X1 U2017 ( .A1(reg_mem[706]), .A2(n3134), .B1(n7026), .B2(data_w[2]), 
        .ZN(n3136) );
  INV_X1 U2018 ( .A(n3137), .ZN(n7021) );
  AOI22_X1 U2019 ( .A1(reg_mem[707]), .A2(n3134), .B1(n7026), .B2(data_w[3]), 
        .ZN(n3137) );
  INV_X1 U2020 ( .A(n3138), .ZN(n7022) );
  AOI22_X1 U2021 ( .A1(reg_mem[708]), .A2(n3134), .B1(n7026), .B2(data_w[4]), 
        .ZN(n3138) );
  INV_X1 U2022 ( .A(n3139), .ZN(n7023) );
  AOI22_X1 U2023 ( .A1(reg_mem[709]), .A2(n3134), .B1(n7026), .B2(data_w[5]), 
        .ZN(n3139) );
  INV_X1 U2024 ( .A(n3140), .ZN(n7024) );
  AOI22_X1 U2025 ( .A1(reg_mem[710]), .A2(n3134), .B1(n7026), .B2(data_w[6]), 
        .ZN(n3140) );
  INV_X1 U2026 ( .A(n3141), .ZN(n7025) );
  AOI22_X1 U2027 ( .A1(reg_mem[711]), .A2(n3134), .B1(n7026), .B2(data_w[7]), 
        .ZN(n3141) );
  INV_X1 U2028 ( .A(n3142), .ZN(n8747) );
  AOI22_X1 U2029 ( .A1(reg_mem[712]), .A2(n3143), .B1(n8755), .B2(data_w[0]), 
        .ZN(n3142) );
  INV_X1 U2030 ( .A(n3144), .ZN(n8748) );
  AOI22_X1 U2031 ( .A1(reg_mem[713]), .A2(n3143), .B1(n8755), .B2(data_w[1]), 
        .ZN(n3144) );
  INV_X1 U2032 ( .A(n3145), .ZN(n8749) );
  AOI22_X1 U2033 ( .A1(reg_mem[714]), .A2(n3143), .B1(n8755), .B2(data_w[2]), 
        .ZN(n3145) );
  INV_X1 U2034 ( .A(n3146), .ZN(n8750) );
  AOI22_X1 U2035 ( .A1(reg_mem[715]), .A2(n3143), .B1(n8755), .B2(data_w[3]), 
        .ZN(n3146) );
  INV_X1 U2036 ( .A(n3147), .ZN(n8751) );
  AOI22_X1 U2037 ( .A1(reg_mem[716]), .A2(n3143), .B1(n8755), .B2(data_w[4]), 
        .ZN(n3147) );
  INV_X1 U2038 ( .A(n3148), .ZN(n8752) );
  AOI22_X1 U2039 ( .A1(reg_mem[717]), .A2(n3143), .B1(n8755), .B2(data_w[5]), 
        .ZN(n3148) );
  INV_X1 U2040 ( .A(n3149), .ZN(n8753) );
  AOI22_X1 U2041 ( .A1(reg_mem[718]), .A2(n3143), .B1(n8755), .B2(data_w[6]), 
        .ZN(n3149) );
  INV_X1 U2042 ( .A(n3150), .ZN(n8754) );
  AOI22_X1 U2043 ( .A1(reg_mem[719]), .A2(n3143), .B1(n8755), .B2(data_w[7]), 
        .ZN(n3150) );
  INV_X1 U2044 ( .A(n3151), .ZN(n7594) );
  AOI22_X1 U2045 ( .A1(reg_mem[720]), .A2(n3152), .B1(n7602), .B2(data_w[0]), 
        .ZN(n3151) );
  INV_X1 U2046 ( .A(n3153), .ZN(n7595) );
  AOI22_X1 U2047 ( .A1(reg_mem[721]), .A2(n3152), .B1(n7602), .B2(data_w[1]), 
        .ZN(n3153) );
  INV_X1 U2048 ( .A(n3154), .ZN(n7596) );
  AOI22_X1 U2049 ( .A1(reg_mem[722]), .A2(n3152), .B1(n7602), .B2(data_w[2]), 
        .ZN(n3154) );
  INV_X1 U2050 ( .A(n3155), .ZN(n7597) );
  AOI22_X1 U2051 ( .A1(reg_mem[723]), .A2(n3152), .B1(n7602), .B2(data_w[3]), 
        .ZN(n3155) );
  INV_X1 U2052 ( .A(n3156), .ZN(n7598) );
  AOI22_X1 U2053 ( .A1(reg_mem[724]), .A2(n3152), .B1(n7602), .B2(data_w[4]), 
        .ZN(n3156) );
  INV_X1 U2054 ( .A(n3157), .ZN(n7599) );
  AOI22_X1 U2055 ( .A1(reg_mem[725]), .A2(n3152), .B1(n7602), .B2(data_w[5]), 
        .ZN(n3157) );
  INV_X1 U2056 ( .A(n3158), .ZN(n7600) );
  AOI22_X1 U2057 ( .A1(reg_mem[726]), .A2(n3152), .B1(n7602), .B2(data_w[6]), 
        .ZN(n3158) );
  INV_X1 U2058 ( .A(n3159), .ZN(n7601) );
  AOI22_X1 U2059 ( .A1(reg_mem[727]), .A2(n3152), .B1(n7602), .B2(data_w[7]), 
        .ZN(n3159) );
  INV_X1 U2060 ( .A(n3160), .ZN(n8171) );
  AOI22_X1 U2061 ( .A1(reg_mem[728]), .A2(n3161), .B1(n8179), .B2(data_w[0]), 
        .ZN(n3160) );
  INV_X1 U2062 ( .A(n3162), .ZN(n8172) );
  AOI22_X1 U2063 ( .A1(reg_mem[729]), .A2(n3161), .B1(n8179), .B2(data_w[1]), 
        .ZN(n3162) );
  INV_X1 U2064 ( .A(n3163), .ZN(n8173) );
  AOI22_X1 U2065 ( .A1(reg_mem[730]), .A2(n3161), .B1(n8179), .B2(data_w[2]), 
        .ZN(n3163) );
  INV_X1 U2066 ( .A(n3164), .ZN(n8174) );
  AOI22_X1 U2067 ( .A1(reg_mem[731]), .A2(n3161), .B1(n8179), .B2(data_w[3]), 
        .ZN(n3164) );
  INV_X1 U2068 ( .A(n3165), .ZN(n8175) );
  AOI22_X1 U2069 ( .A1(reg_mem[732]), .A2(n3161), .B1(n8179), .B2(data_w[4]), 
        .ZN(n3165) );
  INV_X1 U2070 ( .A(n3166), .ZN(n8176) );
  AOI22_X1 U2071 ( .A1(reg_mem[733]), .A2(n3161), .B1(n8179), .B2(data_w[5]), 
        .ZN(n3166) );
  INV_X1 U2072 ( .A(n3167), .ZN(n8177) );
  AOI22_X1 U2073 ( .A1(reg_mem[734]), .A2(n3161), .B1(n8179), .B2(data_w[6]), 
        .ZN(n3167) );
  INV_X1 U2074 ( .A(n3168), .ZN(n8178) );
  AOI22_X1 U2075 ( .A1(reg_mem[735]), .A2(n3161), .B1(n8179), .B2(data_w[7]), 
        .ZN(n3168) );
  INV_X1 U2076 ( .A(n3169), .ZN(n6874) );
  AOI22_X1 U2077 ( .A1(reg_mem[736]), .A2(n3170), .B1(n6882), .B2(data_w[0]), 
        .ZN(n3169) );
  INV_X1 U2078 ( .A(n3171), .ZN(n6875) );
  AOI22_X1 U2079 ( .A1(reg_mem[737]), .A2(n3170), .B1(n6882), .B2(data_w[1]), 
        .ZN(n3171) );
  INV_X1 U2080 ( .A(n3172), .ZN(n6876) );
  AOI22_X1 U2081 ( .A1(reg_mem[738]), .A2(n3170), .B1(n6882), .B2(data_w[2]), 
        .ZN(n3172) );
  INV_X1 U2082 ( .A(n3173), .ZN(n6877) );
  AOI22_X1 U2083 ( .A1(reg_mem[739]), .A2(n3170), .B1(n6882), .B2(data_w[3]), 
        .ZN(n3173) );
  INV_X1 U2084 ( .A(n3174), .ZN(n6878) );
  AOI22_X1 U2085 ( .A1(reg_mem[740]), .A2(n3170), .B1(n6882), .B2(data_w[4]), 
        .ZN(n3174) );
  INV_X1 U2086 ( .A(n3175), .ZN(n6879) );
  AOI22_X1 U2087 ( .A1(reg_mem[741]), .A2(n3170), .B1(n6882), .B2(data_w[5]), 
        .ZN(n3175) );
  INV_X1 U2088 ( .A(n3176), .ZN(n6880) );
  AOI22_X1 U2089 ( .A1(reg_mem[742]), .A2(n3170), .B1(n6882), .B2(data_w[6]), 
        .ZN(n3176) );
  INV_X1 U2090 ( .A(n3177), .ZN(n6881) );
  AOI22_X1 U2091 ( .A1(reg_mem[743]), .A2(n3170), .B1(n6882), .B2(data_w[7]), 
        .ZN(n3177) );
  INV_X1 U2092 ( .A(n3178), .ZN(n8603) );
  AOI22_X1 U2093 ( .A1(reg_mem[744]), .A2(n3179), .B1(n8611), .B2(data_w[0]), 
        .ZN(n3178) );
  INV_X1 U2094 ( .A(n3180), .ZN(n8604) );
  AOI22_X1 U2095 ( .A1(reg_mem[745]), .A2(n3179), .B1(n8611), .B2(data_w[1]), 
        .ZN(n3180) );
  INV_X1 U2096 ( .A(n3181), .ZN(n8605) );
  AOI22_X1 U2097 ( .A1(reg_mem[746]), .A2(n3179), .B1(n8611), .B2(data_w[2]), 
        .ZN(n3181) );
  INV_X1 U2098 ( .A(n3182), .ZN(n8606) );
  AOI22_X1 U2099 ( .A1(reg_mem[747]), .A2(n3179), .B1(n8611), .B2(data_w[3]), 
        .ZN(n3182) );
  INV_X1 U2100 ( .A(n3183), .ZN(n8607) );
  AOI22_X1 U2101 ( .A1(reg_mem[748]), .A2(n3179), .B1(n8611), .B2(data_w[4]), 
        .ZN(n3183) );
  INV_X1 U2102 ( .A(n3184), .ZN(n8608) );
  AOI22_X1 U2103 ( .A1(reg_mem[749]), .A2(n3179), .B1(n8611), .B2(data_w[5]), 
        .ZN(n3184) );
  INV_X1 U2104 ( .A(n3185), .ZN(n8609) );
  AOI22_X1 U2105 ( .A1(reg_mem[750]), .A2(n3179), .B1(n8611), .B2(data_w[6]), 
        .ZN(n3185) );
  INV_X1 U2106 ( .A(n3186), .ZN(n8610) );
  AOI22_X1 U2107 ( .A1(reg_mem[751]), .A2(n3179), .B1(n8611), .B2(data_w[7]), 
        .ZN(n3186) );
  INV_X1 U2108 ( .A(n3187), .ZN(n7450) );
  AOI22_X1 U2109 ( .A1(reg_mem[752]), .A2(n3188), .B1(n7458), .B2(data_w[0]), 
        .ZN(n3187) );
  INV_X1 U2110 ( .A(n3189), .ZN(n7451) );
  AOI22_X1 U2111 ( .A1(reg_mem[753]), .A2(n3188), .B1(n7458), .B2(data_w[1]), 
        .ZN(n3189) );
  INV_X1 U2112 ( .A(n3190), .ZN(n7452) );
  AOI22_X1 U2113 ( .A1(reg_mem[754]), .A2(n3188), .B1(n7458), .B2(data_w[2]), 
        .ZN(n3190) );
  INV_X1 U2114 ( .A(n3191), .ZN(n7453) );
  AOI22_X1 U2115 ( .A1(reg_mem[755]), .A2(n3188), .B1(n7458), .B2(data_w[3]), 
        .ZN(n3191) );
  INV_X1 U2116 ( .A(n3192), .ZN(n7454) );
  AOI22_X1 U2117 ( .A1(reg_mem[756]), .A2(n3188), .B1(n7458), .B2(data_w[4]), 
        .ZN(n3192) );
  INV_X1 U2118 ( .A(n3193), .ZN(n7455) );
  AOI22_X1 U2119 ( .A1(reg_mem[757]), .A2(n3188), .B1(n7458), .B2(data_w[5]), 
        .ZN(n3193) );
  INV_X1 U2120 ( .A(n3194), .ZN(n7456) );
  AOI22_X1 U2121 ( .A1(reg_mem[758]), .A2(n3188), .B1(n7458), .B2(data_w[6]), 
        .ZN(n3194) );
  INV_X1 U2122 ( .A(n3195), .ZN(n7457) );
  AOI22_X1 U2123 ( .A1(reg_mem[759]), .A2(n3188), .B1(n7458), .B2(data_w[7]), 
        .ZN(n3195) );
  INV_X1 U2124 ( .A(n3196), .ZN(n8027) );
  AOI22_X1 U2125 ( .A1(reg_mem[760]), .A2(n3197), .B1(n8035), .B2(data_w[0]), 
        .ZN(n3196) );
  INV_X1 U2126 ( .A(n3198), .ZN(n8028) );
  AOI22_X1 U2127 ( .A1(reg_mem[761]), .A2(n3197), .B1(n8035), .B2(data_w[1]), 
        .ZN(n3198) );
  INV_X1 U2128 ( .A(n3199), .ZN(n8029) );
  AOI22_X1 U2129 ( .A1(reg_mem[762]), .A2(n3197), .B1(n8035), .B2(data_w[2]), 
        .ZN(n3199) );
  INV_X1 U2130 ( .A(n3200), .ZN(n8030) );
  AOI22_X1 U2131 ( .A1(reg_mem[763]), .A2(n3197), .B1(n8035), .B2(data_w[3]), 
        .ZN(n3200) );
  INV_X1 U2132 ( .A(n3201), .ZN(n8031) );
  AOI22_X1 U2133 ( .A1(reg_mem[764]), .A2(n3197), .B1(n8035), .B2(data_w[4]), 
        .ZN(n3201) );
  INV_X1 U2134 ( .A(n3202), .ZN(n8032) );
  AOI22_X1 U2135 ( .A1(reg_mem[765]), .A2(n3197), .B1(n8035), .B2(data_w[5]), 
        .ZN(n3202) );
  INV_X1 U2136 ( .A(n3203), .ZN(n8033) );
  AOI22_X1 U2137 ( .A1(reg_mem[766]), .A2(n3197), .B1(n8035), .B2(data_w[6]), 
        .ZN(n3203) );
  INV_X1 U2138 ( .A(n3204), .ZN(n8034) );
  AOI22_X1 U2139 ( .A1(reg_mem[767]), .A2(n3197), .B1(n8035), .B2(data_w[7]), 
        .ZN(n3204) );
  INV_X1 U2140 ( .A(n3205), .ZN(n7297) );
  AOI22_X1 U2141 ( .A1(reg_mem[768]), .A2(n3206), .B1(n7305), .B2(data_w[0]), 
        .ZN(n3205) );
  INV_X1 U2142 ( .A(n3207), .ZN(n7298) );
  AOI22_X1 U2143 ( .A1(reg_mem[769]), .A2(n3206), .B1(n7305), .B2(data_w[1]), 
        .ZN(n3207) );
  INV_X1 U2144 ( .A(n3208), .ZN(n7299) );
  AOI22_X1 U2145 ( .A1(reg_mem[770]), .A2(n3206), .B1(n7305), .B2(data_w[2]), 
        .ZN(n3208) );
  INV_X1 U2146 ( .A(n3209), .ZN(n7300) );
  AOI22_X1 U2147 ( .A1(reg_mem[771]), .A2(n3206), .B1(n7305), .B2(data_w[3]), 
        .ZN(n3209) );
  INV_X1 U2148 ( .A(n3210), .ZN(n7301) );
  AOI22_X1 U2149 ( .A1(reg_mem[772]), .A2(n3206), .B1(n7305), .B2(data_w[4]), 
        .ZN(n3210) );
  INV_X1 U2150 ( .A(n3211), .ZN(n7302) );
  AOI22_X1 U2151 ( .A1(reg_mem[773]), .A2(n3206), .B1(n7305), .B2(data_w[5]), 
        .ZN(n3211) );
  INV_X1 U2152 ( .A(n3212), .ZN(n7303) );
  AOI22_X1 U2153 ( .A1(reg_mem[774]), .A2(n3206), .B1(n7305), .B2(data_w[6]), 
        .ZN(n3212) );
  INV_X1 U2154 ( .A(n3213), .ZN(n7304) );
  AOI22_X1 U2155 ( .A1(reg_mem[775]), .A2(n3206), .B1(n7305), .B2(data_w[7]), 
        .ZN(n3213) );
  INV_X1 U2156 ( .A(n3215), .ZN(n9026) );
  AOI22_X1 U2157 ( .A1(reg_mem[776]), .A2(n3216), .B1(n9034), .B2(data_w[0]), 
        .ZN(n3215) );
  INV_X1 U2158 ( .A(n3217), .ZN(n9027) );
  AOI22_X1 U2159 ( .A1(reg_mem[777]), .A2(n3216), .B1(n9034), .B2(data_w[1]), 
        .ZN(n3217) );
  INV_X1 U2160 ( .A(n3218), .ZN(n9028) );
  AOI22_X1 U2161 ( .A1(reg_mem[778]), .A2(n3216), .B1(n9034), .B2(data_w[2]), 
        .ZN(n3218) );
  INV_X1 U2162 ( .A(n3219), .ZN(n9029) );
  AOI22_X1 U2163 ( .A1(reg_mem[779]), .A2(n3216), .B1(n9034), .B2(data_w[3]), 
        .ZN(n3219) );
  INV_X1 U2164 ( .A(n3220), .ZN(n9030) );
  AOI22_X1 U2165 ( .A1(reg_mem[780]), .A2(n3216), .B1(n9034), .B2(data_w[4]), 
        .ZN(n3220) );
  INV_X1 U2166 ( .A(n3221), .ZN(n9031) );
  AOI22_X1 U2167 ( .A1(reg_mem[781]), .A2(n3216), .B1(n9034), .B2(data_w[5]), 
        .ZN(n3221) );
  INV_X1 U2168 ( .A(n3222), .ZN(n9032) );
  AOI22_X1 U2169 ( .A1(reg_mem[782]), .A2(n3216), .B1(n9034), .B2(data_w[6]), 
        .ZN(n3222) );
  INV_X1 U2170 ( .A(n3223), .ZN(n9033) );
  AOI22_X1 U2171 ( .A1(reg_mem[783]), .A2(n3216), .B1(n9034), .B2(data_w[7]), 
        .ZN(n3223) );
  INV_X1 U2172 ( .A(n3224), .ZN(n7873) );
  AOI22_X1 U2173 ( .A1(reg_mem[784]), .A2(n3225), .B1(n7881), .B2(data_w[0]), 
        .ZN(n3224) );
  INV_X1 U2174 ( .A(n3226), .ZN(n7874) );
  AOI22_X1 U2175 ( .A1(reg_mem[785]), .A2(n3225), .B1(n7881), .B2(data_w[1]), 
        .ZN(n3226) );
  INV_X1 U2176 ( .A(n3227), .ZN(n7875) );
  AOI22_X1 U2177 ( .A1(reg_mem[786]), .A2(n3225), .B1(n7881), .B2(data_w[2]), 
        .ZN(n3227) );
  INV_X1 U2178 ( .A(n3228), .ZN(n7876) );
  AOI22_X1 U2179 ( .A1(reg_mem[787]), .A2(n3225), .B1(n7881), .B2(data_w[3]), 
        .ZN(n3228) );
  INV_X1 U2180 ( .A(n3229), .ZN(n7877) );
  AOI22_X1 U2181 ( .A1(reg_mem[788]), .A2(n3225), .B1(n7881), .B2(data_w[4]), 
        .ZN(n3229) );
  INV_X1 U2182 ( .A(n3230), .ZN(n7878) );
  AOI22_X1 U2183 ( .A1(reg_mem[789]), .A2(n3225), .B1(n7881), .B2(data_w[5]), 
        .ZN(n3230) );
  INV_X1 U2184 ( .A(n3231), .ZN(n7879) );
  AOI22_X1 U2185 ( .A1(reg_mem[790]), .A2(n3225), .B1(n7881), .B2(data_w[6]), 
        .ZN(n3231) );
  INV_X1 U2186 ( .A(n3232), .ZN(n7880) );
  AOI22_X1 U2187 ( .A1(reg_mem[791]), .A2(n3225), .B1(n7881), .B2(data_w[7]), 
        .ZN(n3232) );
  INV_X1 U2188 ( .A(n3233), .ZN(n8450) );
  AOI22_X1 U2189 ( .A1(reg_mem[792]), .A2(n3234), .B1(n8458), .B2(data_w[0]), 
        .ZN(n3233) );
  INV_X1 U2190 ( .A(n3235), .ZN(n8451) );
  AOI22_X1 U2191 ( .A1(reg_mem[793]), .A2(n3234), .B1(n8458), .B2(data_w[1]), 
        .ZN(n3235) );
  INV_X1 U2192 ( .A(n3236), .ZN(n8452) );
  AOI22_X1 U2193 ( .A1(reg_mem[794]), .A2(n3234), .B1(n8458), .B2(data_w[2]), 
        .ZN(n3236) );
  INV_X1 U2194 ( .A(n3237), .ZN(n8453) );
  AOI22_X1 U2195 ( .A1(reg_mem[795]), .A2(n3234), .B1(n8458), .B2(data_w[3]), 
        .ZN(n3237) );
  INV_X1 U2196 ( .A(n3238), .ZN(n8454) );
  AOI22_X1 U2197 ( .A1(reg_mem[796]), .A2(n3234), .B1(n8458), .B2(data_w[4]), 
        .ZN(n3238) );
  INV_X1 U2198 ( .A(n3239), .ZN(n8455) );
  AOI22_X1 U2199 ( .A1(reg_mem[797]), .A2(n3234), .B1(n8458), .B2(data_w[5]), 
        .ZN(n3239) );
  INV_X1 U2200 ( .A(n3240), .ZN(n8456) );
  AOI22_X1 U2201 ( .A1(reg_mem[798]), .A2(n3234), .B1(n8458), .B2(data_w[6]), 
        .ZN(n3240) );
  INV_X1 U2202 ( .A(n3241), .ZN(n8457) );
  AOI22_X1 U2203 ( .A1(reg_mem[799]), .A2(n3234), .B1(n8458), .B2(data_w[7]), 
        .ZN(n3241) );
  INV_X1 U2204 ( .A(n3242), .ZN(n7153) );
  AOI22_X1 U2205 ( .A1(reg_mem[800]), .A2(n3243), .B1(n7161), .B2(data_w[0]), 
        .ZN(n3242) );
  INV_X1 U2206 ( .A(n3244), .ZN(n7154) );
  AOI22_X1 U2207 ( .A1(reg_mem[801]), .A2(n3243), .B1(n7161), .B2(data_w[1]), 
        .ZN(n3244) );
  INV_X1 U2208 ( .A(n3245), .ZN(n7155) );
  AOI22_X1 U2209 ( .A1(reg_mem[802]), .A2(n3243), .B1(n7161), .B2(data_w[2]), 
        .ZN(n3245) );
  INV_X1 U2210 ( .A(n3246), .ZN(n7156) );
  AOI22_X1 U2211 ( .A1(reg_mem[803]), .A2(n3243), .B1(n7161), .B2(data_w[3]), 
        .ZN(n3246) );
  INV_X1 U2212 ( .A(n3247), .ZN(n7157) );
  AOI22_X1 U2213 ( .A1(reg_mem[804]), .A2(n3243), .B1(n7161), .B2(data_w[4]), 
        .ZN(n3247) );
  INV_X1 U2214 ( .A(n3248), .ZN(n7158) );
  AOI22_X1 U2215 ( .A1(reg_mem[805]), .A2(n3243), .B1(n7161), .B2(data_w[5]), 
        .ZN(n3248) );
  INV_X1 U2216 ( .A(n3249), .ZN(n7159) );
  AOI22_X1 U2217 ( .A1(reg_mem[806]), .A2(n3243), .B1(n7161), .B2(data_w[6]), 
        .ZN(n3249) );
  INV_X1 U2218 ( .A(n3250), .ZN(n7160) );
  AOI22_X1 U2219 ( .A1(reg_mem[807]), .A2(n3243), .B1(n7161), .B2(data_w[7]), 
        .ZN(n3250) );
  INV_X1 U2220 ( .A(n3251), .ZN(n8882) );
  AOI22_X1 U2221 ( .A1(reg_mem[808]), .A2(n3252), .B1(n8890), .B2(data_w[0]), 
        .ZN(n3251) );
  INV_X1 U2222 ( .A(n3253), .ZN(n8883) );
  AOI22_X1 U2223 ( .A1(reg_mem[809]), .A2(n3252), .B1(n8890), .B2(data_w[1]), 
        .ZN(n3253) );
  INV_X1 U2224 ( .A(n3254), .ZN(n8884) );
  AOI22_X1 U2225 ( .A1(reg_mem[810]), .A2(n3252), .B1(n8890), .B2(data_w[2]), 
        .ZN(n3254) );
  INV_X1 U2226 ( .A(n3255), .ZN(n8885) );
  AOI22_X1 U2227 ( .A1(reg_mem[811]), .A2(n3252), .B1(n8890), .B2(data_w[3]), 
        .ZN(n3255) );
  INV_X1 U2228 ( .A(n3256), .ZN(n8886) );
  AOI22_X1 U2229 ( .A1(reg_mem[812]), .A2(n3252), .B1(n8890), .B2(data_w[4]), 
        .ZN(n3256) );
  INV_X1 U2230 ( .A(n3257), .ZN(n8887) );
  AOI22_X1 U2231 ( .A1(reg_mem[813]), .A2(n3252), .B1(n8890), .B2(data_w[5]), 
        .ZN(n3257) );
  INV_X1 U2232 ( .A(n3258), .ZN(n8888) );
  AOI22_X1 U2233 ( .A1(reg_mem[814]), .A2(n3252), .B1(n8890), .B2(data_w[6]), 
        .ZN(n3258) );
  INV_X1 U2234 ( .A(n3259), .ZN(n8889) );
  AOI22_X1 U2235 ( .A1(reg_mem[815]), .A2(n3252), .B1(n8890), .B2(data_w[7]), 
        .ZN(n3259) );
  INV_X1 U2236 ( .A(n3260), .ZN(n7729) );
  AOI22_X1 U2237 ( .A1(reg_mem[816]), .A2(n3261), .B1(n7737), .B2(data_w[0]), 
        .ZN(n3260) );
  INV_X1 U2238 ( .A(n3262), .ZN(n7730) );
  AOI22_X1 U2239 ( .A1(reg_mem[817]), .A2(n3261), .B1(n7737), .B2(data_w[1]), 
        .ZN(n3262) );
  INV_X1 U2240 ( .A(n3263), .ZN(n7731) );
  AOI22_X1 U2241 ( .A1(reg_mem[818]), .A2(n3261), .B1(n7737), .B2(data_w[2]), 
        .ZN(n3263) );
  INV_X1 U2242 ( .A(n3264), .ZN(n7732) );
  AOI22_X1 U2243 ( .A1(reg_mem[819]), .A2(n3261), .B1(n7737), .B2(data_w[3]), 
        .ZN(n3264) );
  INV_X1 U2244 ( .A(n3265), .ZN(n7733) );
  AOI22_X1 U2245 ( .A1(reg_mem[820]), .A2(n3261), .B1(n7737), .B2(data_w[4]), 
        .ZN(n3265) );
  INV_X1 U2246 ( .A(n3266), .ZN(n7734) );
  AOI22_X1 U2247 ( .A1(reg_mem[821]), .A2(n3261), .B1(n7737), .B2(data_w[5]), 
        .ZN(n3266) );
  INV_X1 U2248 ( .A(n3267), .ZN(n7735) );
  AOI22_X1 U2249 ( .A1(reg_mem[822]), .A2(n3261), .B1(n7737), .B2(data_w[6]), 
        .ZN(n3267) );
  INV_X1 U2250 ( .A(n3268), .ZN(n7736) );
  AOI22_X1 U2251 ( .A1(reg_mem[823]), .A2(n3261), .B1(n7737), .B2(data_w[7]), 
        .ZN(n3268) );
  INV_X1 U2252 ( .A(n3269), .ZN(n8306) );
  AOI22_X1 U2253 ( .A1(reg_mem[824]), .A2(n3270), .B1(n8314), .B2(data_w[0]), 
        .ZN(n3269) );
  INV_X1 U2254 ( .A(n3271), .ZN(n8307) );
  AOI22_X1 U2255 ( .A1(reg_mem[825]), .A2(n3270), .B1(n8314), .B2(data_w[1]), 
        .ZN(n3271) );
  INV_X1 U2256 ( .A(n3272), .ZN(n8308) );
  AOI22_X1 U2257 ( .A1(reg_mem[826]), .A2(n3270), .B1(n8314), .B2(data_w[2]), 
        .ZN(n3272) );
  INV_X1 U2258 ( .A(n3273), .ZN(n8309) );
  AOI22_X1 U2259 ( .A1(reg_mem[827]), .A2(n3270), .B1(n8314), .B2(data_w[3]), 
        .ZN(n3273) );
  INV_X1 U2260 ( .A(n3274), .ZN(n8310) );
  AOI22_X1 U2261 ( .A1(reg_mem[828]), .A2(n3270), .B1(n8314), .B2(data_w[4]), 
        .ZN(n3274) );
  INV_X1 U2262 ( .A(n3275), .ZN(n8311) );
  AOI22_X1 U2263 ( .A1(reg_mem[829]), .A2(n3270), .B1(n8314), .B2(data_w[5]), 
        .ZN(n3275) );
  INV_X1 U2264 ( .A(n3276), .ZN(n8312) );
  AOI22_X1 U2265 ( .A1(reg_mem[830]), .A2(n3270), .B1(n8314), .B2(data_w[6]), 
        .ZN(n3276) );
  INV_X1 U2266 ( .A(n3277), .ZN(n8313) );
  AOI22_X1 U2267 ( .A1(reg_mem[831]), .A2(n3270), .B1(n8314), .B2(data_w[7]), 
        .ZN(n3277) );
  INV_X1 U2268 ( .A(n3278), .ZN(n7009) );
  AOI22_X1 U2269 ( .A1(reg_mem[832]), .A2(n3279), .B1(n7017), .B2(data_w[0]), 
        .ZN(n3278) );
  INV_X1 U2270 ( .A(n3280), .ZN(n7010) );
  AOI22_X1 U2271 ( .A1(reg_mem[833]), .A2(n3279), .B1(n7017), .B2(data_w[1]), 
        .ZN(n3280) );
  INV_X1 U2272 ( .A(n3281), .ZN(n7011) );
  AOI22_X1 U2273 ( .A1(reg_mem[834]), .A2(n3279), .B1(n7017), .B2(data_w[2]), 
        .ZN(n3281) );
  INV_X1 U2274 ( .A(n3282), .ZN(n7012) );
  AOI22_X1 U2275 ( .A1(reg_mem[835]), .A2(n3279), .B1(n7017), .B2(data_w[3]), 
        .ZN(n3282) );
  INV_X1 U2276 ( .A(n3283), .ZN(n7013) );
  AOI22_X1 U2277 ( .A1(reg_mem[836]), .A2(n3279), .B1(n7017), .B2(data_w[4]), 
        .ZN(n3283) );
  INV_X1 U2278 ( .A(n3284), .ZN(n7014) );
  AOI22_X1 U2279 ( .A1(reg_mem[837]), .A2(n3279), .B1(n7017), .B2(data_w[5]), 
        .ZN(n3284) );
  INV_X1 U2280 ( .A(n3285), .ZN(n7015) );
  AOI22_X1 U2281 ( .A1(reg_mem[838]), .A2(n3279), .B1(n7017), .B2(data_w[6]), 
        .ZN(n3285) );
  INV_X1 U2282 ( .A(n3286), .ZN(n7016) );
  AOI22_X1 U2283 ( .A1(reg_mem[839]), .A2(n3279), .B1(n7017), .B2(data_w[7]), 
        .ZN(n3286) );
  INV_X1 U2284 ( .A(n3287), .ZN(n8738) );
  AOI22_X1 U2285 ( .A1(reg_mem[840]), .A2(n3288), .B1(n8746), .B2(data_w[0]), 
        .ZN(n3287) );
  INV_X1 U2286 ( .A(n3289), .ZN(n8739) );
  AOI22_X1 U2287 ( .A1(reg_mem[841]), .A2(n3288), .B1(n8746), .B2(data_w[1]), 
        .ZN(n3289) );
  INV_X1 U2288 ( .A(n3290), .ZN(n8740) );
  AOI22_X1 U2289 ( .A1(reg_mem[842]), .A2(n3288), .B1(n8746), .B2(data_w[2]), 
        .ZN(n3290) );
  INV_X1 U2290 ( .A(n3291), .ZN(n8741) );
  AOI22_X1 U2291 ( .A1(reg_mem[843]), .A2(n3288), .B1(n8746), .B2(data_w[3]), 
        .ZN(n3291) );
  INV_X1 U2292 ( .A(n3292), .ZN(n8742) );
  AOI22_X1 U2293 ( .A1(reg_mem[844]), .A2(n3288), .B1(n8746), .B2(data_w[4]), 
        .ZN(n3292) );
  INV_X1 U2294 ( .A(n3293), .ZN(n8743) );
  AOI22_X1 U2295 ( .A1(reg_mem[845]), .A2(n3288), .B1(n8746), .B2(data_w[5]), 
        .ZN(n3293) );
  INV_X1 U2296 ( .A(n3294), .ZN(n8744) );
  AOI22_X1 U2297 ( .A1(reg_mem[846]), .A2(n3288), .B1(n8746), .B2(data_w[6]), 
        .ZN(n3294) );
  INV_X1 U2298 ( .A(n3295), .ZN(n8745) );
  AOI22_X1 U2299 ( .A1(reg_mem[847]), .A2(n3288), .B1(n8746), .B2(data_w[7]), 
        .ZN(n3295) );
  INV_X1 U2300 ( .A(n3296), .ZN(n7585) );
  AOI22_X1 U2301 ( .A1(reg_mem[848]), .A2(n3297), .B1(n7593), .B2(data_w[0]), 
        .ZN(n3296) );
  INV_X1 U2302 ( .A(n3298), .ZN(n7586) );
  AOI22_X1 U2303 ( .A1(reg_mem[849]), .A2(n3297), .B1(n7593), .B2(data_w[1]), 
        .ZN(n3298) );
  INV_X1 U2304 ( .A(n3299), .ZN(n7587) );
  AOI22_X1 U2305 ( .A1(reg_mem[850]), .A2(n3297), .B1(n7593), .B2(data_w[2]), 
        .ZN(n3299) );
  INV_X1 U2306 ( .A(n3300), .ZN(n7588) );
  AOI22_X1 U2307 ( .A1(reg_mem[851]), .A2(n3297), .B1(n7593), .B2(data_w[3]), 
        .ZN(n3300) );
  INV_X1 U2308 ( .A(n3301), .ZN(n7589) );
  AOI22_X1 U2309 ( .A1(reg_mem[852]), .A2(n3297), .B1(n7593), .B2(data_w[4]), 
        .ZN(n3301) );
  INV_X1 U2310 ( .A(n3302), .ZN(n7590) );
  AOI22_X1 U2311 ( .A1(reg_mem[853]), .A2(n3297), .B1(n7593), .B2(data_w[5]), 
        .ZN(n3302) );
  INV_X1 U2312 ( .A(n3303), .ZN(n7591) );
  AOI22_X1 U2313 ( .A1(reg_mem[854]), .A2(n3297), .B1(n7593), .B2(data_w[6]), 
        .ZN(n3303) );
  INV_X1 U2314 ( .A(n3304), .ZN(n7592) );
  AOI22_X1 U2315 ( .A1(reg_mem[855]), .A2(n3297), .B1(n7593), .B2(data_w[7]), 
        .ZN(n3304) );
  INV_X1 U2316 ( .A(n3305), .ZN(n8162) );
  AOI22_X1 U2317 ( .A1(reg_mem[856]), .A2(n3306), .B1(n8170), .B2(data_w[0]), 
        .ZN(n3305) );
  INV_X1 U2318 ( .A(n3307), .ZN(n8163) );
  AOI22_X1 U2319 ( .A1(reg_mem[857]), .A2(n3306), .B1(n8170), .B2(data_w[1]), 
        .ZN(n3307) );
  INV_X1 U2320 ( .A(n3308), .ZN(n8164) );
  AOI22_X1 U2321 ( .A1(reg_mem[858]), .A2(n3306), .B1(n8170), .B2(data_w[2]), 
        .ZN(n3308) );
  INV_X1 U2322 ( .A(n3309), .ZN(n8165) );
  AOI22_X1 U2323 ( .A1(reg_mem[859]), .A2(n3306), .B1(n8170), .B2(data_w[3]), 
        .ZN(n3309) );
  INV_X1 U2324 ( .A(n3310), .ZN(n8166) );
  AOI22_X1 U2325 ( .A1(reg_mem[860]), .A2(n3306), .B1(n8170), .B2(data_w[4]), 
        .ZN(n3310) );
  INV_X1 U2326 ( .A(n3311), .ZN(n8167) );
  AOI22_X1 U2327 ( .A1(reg_mem[861]), .A2(n3306), .B1(n8170), .B2(data_w[5]), 
        .ZN(n3311) );
  INV_X1 U2328 ( .A(n3312), .ZN(n8168) );
  AOI22_X1 U2329 ( .A1(reg_mem[862]), .A2(n3306), .B1(n8170), .B2(data_w[6]), 
        .ZN(n3312) );
  INV_X1 U2330 ( .A(n3313), .ZN(n8169) );
  AOI22_X1 U2331 ( .A1(reg_mem[863]), .A2(n3306), .B1(n8170), .B2(data_w[7]), 
        .ZN(n3313) );
  INV_X1 U2332 ( .A(n3314), .ZN(n6865) );
  AOI22_X1 U2333 ( .A1(reg_mem[864]), .A2(n3315), .B1(n6873), .B2(data_w[0]), 
        .ZN(n3314) );
  INV_X1 U2334 ( .A(n3316), .ZN(n6866) );
  AOI22_X1 U2335 ( .A1(reg_mem[865]), .A2(n3315), .B1(n6873), .B2(data_w[1]), 
        .ZN(n3316) );
  INV_X1 U2336 ( .A(n3317), .ZN(n6867) );
  AOI22_X1 U2337 ( .A1(reg_mem[866]), .A2(n3315), .B1(n6873), .B2(data_w[2]), 
        .ZN(n3317) );
  INV_X1 U2338 ( .A(n3318), .ZN(n6868) );
  AOI22_X1 U2339 ( .A1(reg_mem[867]), .A2(n3315), .B1(n6873), .B2(data_w[3]), 
        .ZN(n3318) );
  INV_X1 U2340 ( .A(n3319), .ZN(n6869) );
  AOI22_X1 U2341 ( .A1(reg_mem[868]), .A2(n3315), .B1(n6873), .B2(data_w[4]), 
        .ZN(n3319) );
  INV_X1 U2342 ( .A(n3320), .ZN(n6870) );
  AOI22_X1 U2343 ( .A1(reg_mem[869]), .A2(n3315), .B1(n6873), .B2(data_w[5]), 
        .ZN(n3320) );
  INV_X1 U2344 ( .A(n3321), .ZN(n6871) );
  AOI22_X1 U2345 ( .A1(reg_mem[870]), .A2(n3315), .B1(n6873), .B2(data_w[6]), 
        .ZN(n3321) );
  INV_X1 U2346 ( .A(n3322), .ZN(n6872) );
  AOI22_X1 U2347 ( .A1(reg_mem[871]), .A2(n3315), .B1(n6873), .B2(data_w[7]), 
        .ZN(n3322) );
  INV_X1 U2348 ( .A(n3323), .ZN(n8594) );
  AOI22_X1 U2349 ( .A1(reg_mem[872]), .A2(n3324), .B1(n8602), .B2(data_w[0]), 
        .ZN(n3323) );
  INV_X1 U2350 ( .A(n3325), .ZN(n8595) );
  AOI22_X1 U2351 ( .A1(reg_mem[873]), .A2(n3324), .B1(n8602), .B2(data_w[1]), 
        .ZN(n3325) );
  INV_X1 U2352 ( .A(n3326), .ZN(n8596) );
  AOI22_X1 U2353 ( .A1(reg_mem[874]), .A2(n3324), .B1(n8602), .B2(data_w[2]), 
        .ZN(n3326) );
  INV_X1 U2354 ( .A(n3327), .ZN(n8597) );
  AOI22_X1 U2355 ( .A1(reg_mem[875]), .A2(n3324), .B1(n8602), .B2(data_w[3]), 
        .ZN(n3327) );
  INV_X1 U2356 ( .A(n3328), .ZN(n8598) );
  AOI22_X1 U2357 ( .A1(reg_mem[876]), .A2(n3324), .B1(n8602), .B2(data_w[4]), 
        .ZN(n3328) );
  INV_X1 U2358 ( .A(n3329), .ZN(n8599) );
  AOI22_X1 U2359 ( .A1(reg_mem[877]), .A2(n3324), .B1(n8602), .B2(data_w[5]), 
        .ZN(n3329) );
  INV_X1 U2360 ( .A(n3330), .ZN(n8600) );
  AOI22_X1 U2361 ( .A1(reg_mem[878]), .A2(n3324), .B1(n8602), .B2(data_w[6]), 
        .ZN(n3330) );
  INV_X1 U2362 ( .A(n3331), .ZN(n8601) );
  AOI22_X1 U2363 ( .A1(reg_mem[879]), .A2(n3324), .B1(n8602), .B2(data_w[7]), 
        .ZN(n3331) );
  INV_X1 U2364 ( .A(n3332), .ZN(n7441) );
  AOI22_X1 U2365 ( .A1(reg_mem[880]), .A2(n3333), .B1(n7449), .B2(data_w[0]), 
        .ZN(n3332) );
  INV_X1 U2366 ( .A(n3334), .ZN(n7442) );
  AOI22_X1 U2367 ( .A1(reg_mem[881]), .A2(n3333), .B1(n7449), .B2(data_w[1]), 
        .ZN(n3334) );
  INV_X1 U2368 ( .A(n3335), .ZN(n7443) );
  AOI22_X1 U2369 ( .A1(reg_mem[882]), .A2(n3333), .B1(n7449), .B2(data_w[2]), 
        .ZN(n3335) );
  INV_X1 U2370 ( .A(n3336), .ZN(n7444) );
  AOI22_X1 U2371 ( .A1(reg_mem[883]), .A2(n3333), .B1(n7449), .B2(data_w[3]), 
        .ZN(n3336) );
  INV_X1 U2372 ( .A(n3337), .ZN(n7445) );
  AOI22_X1 U2373 ( .A1(reg_mem[884]), .A2(n3333), .B1(n7449), .B2(data_w[4]), 
        .ZN(n3337) );
  INV_X1 U2374 ( .A(n3338), .ZN(n7446) );
  AOI22_X1 U2375 ( .A1(reg_mem[885]), .A2(n3333), .B1(n7449), .B2(data_w[5]), 
        .ZN(n3338) );
  INV_X1 U2376 ( .A(n3339), .ZN(n7447) );
  AOI22_X1 U2377 ( .A1(reg_mem[886]), .A2(n3333), .B1(n7449), .B2(data_w[6]), 
        .ZN(n3339) );
  INV_X1 U2378 ( .A(n3340), .ZN(n7448) );
  AOI22_X1 U2379 ( .A1(reg_mem[887]), .A2(n3333), .B1(n7449), .B2(data_w[7]), 
        .ZN(n3340) );
  INV_X1 U2380 ( .A(n3341), .ZN(n8018) );
  AOI22_X1 U2381 ( .A1(reg_mem[888]), .A2(n3342), .B1(n8026), .B2(data_w[0]), 
        .ZN(n3341) );
  INV_X1 U2382 ( .A(n3343), .ZN(n8019) );
  AOI22_X1 U2383 ( .A1(reg_mem[889]), .A2(n3342), .B1(n8026), .B2(data_w[1]), 
        .ZN(n3343) );
  INV_X1 U2384 ( .A(n3344), .ZN(n8020) );
  AOI22_X1 U2385 ( .A1(reg_mem[890]), .A2(n3342), .B1(n8026), .B2(data_w[2]), 
        .ZN(n3344) );
  INV_X1 U2386 ( .A(n3345), .ZN(n8021) );
  AOI22_X1 U2387 ( .A1(reg_mem[891]), .A2(n3342), .B1(n8026), .B2(data_w[3]), 
        .ZN(n3345) );
  INV_X1 U2388 ( .A(n3346), .ZN(n8022) );
  AOI22_X1 U2389 ( .A1(reg_mem[892]), .A2(n3342), .B1(n8026), .B2(data_w[4]), 
        .ZN(n3346) );
  INV_X1 U2390 ( .A(n3347), .ZN(n8023) );
  AOI22_X1 U2391 ( .A1(reg_mem[893]), .A2(n3342), .B1(n8026), .B2(data_w[5]), 
        .ZN(n3347) );
  INV_X1 U2392 ( .A(n3348), .ZN(n8024) );
  AOI22_X1 U2393 ( .A1(reg_mem[894]), .A2(n3342), .B1(n8026), .B2(data_w[6]), 
        .ZN(n3348) );
  INV_X1 U2394 ( .A(n3349), .ZN(n8025) );
  AOI22_X1 U2395 ( .A1(reg_mem[895]), .A2(n3342), .B1(n8026), .B2(data_w[7]), 
        .ZN(n3349) );
  INV_X1 U2396 ( .A(n3350), .ZN(n7288) );
  AOI22_X1 U2397 ( .A1(reg_mem[896]), .A2(n3351), .B1(n7296), .B2(data_w[0]), 
        .ZN(n3350) );
  INV_X1 U2398 ( .A(n3352), .ZN(n7289) );
  AOI22_X1 U2399 ( .A1(reg_mem[897]), .A2(n3351), .B1(n7296), .B2(data_w[1]), 
        .ZN(n3352) );
  INV_X1 U2400 ( .A(n3353), .ZN(n7290) );
  AOI22_X1 U2401 ( .A1(reg_mem[898]), .A2(n3351), .B1(n7296), .B2(data_w[2]), 
        .ZN(n3353) );
  INV_X1 U2402 ( .A(n3354), .ZN(n7291) );
  AOI22_X1 U2403 ( .A1(reg_mem[899]), .A2(n3351), .B1(n7296), .B2(data_w[3]), 
        .ZN(n3354) );
  INV_X1 U2404 ( .A(n3355), .ZN(n7292) );
  AOI22_X1 U2405 ( .A1(reg_mem[900]), .A2(n3351), .B1(n7296), .B2(data_w[4]), 
        .ZN(n3355) );
  INV_X1 U2406 ( .A(n3356), .ZN(n7293) );
  AOI22_X1 U2407 ( .A1(reg_mem[901]), .A2(n3351), .B1(n7296), .B2(data_w[5]), 
        .ZN(n3356) );
  INV_X1 U2408 ( .A(n3357), .ZN(n7294) );
  AOI22_X1 U2409 ( .A1(reg_mem[902]), .A2(n3351), .B1(n7296), .B2(data_w[6]), 
        .ZN(n3357) );
  INV_X1 U2410 ( .A(n3358), .ZN(n7295) );
  AOI22_X1 U2411 ( .A1(reg_mem[903]), .A2(n3351), .B1(n7296), .B2(data_w[7]), 
        .ZN(n3358) );
  INV_X1 U2412 ( .A(n3360), .ZN(n9017) );
  AOI22_X1 U2413 ( .A1(reg_mem[904]), .A2(n3361), .B1(n9025), .B2(data_w[0]), 
        .ZN(n3360) );
  INV_X1 U2414 ( .A(n3362), .ZN(n9018) );
  AOI22_X1 U2415 ( .A1(reg_mem[905]), .A2(n3361), .B1(n9025), .B2(data_w[1]), 
        .ZN(n3362) );
  INV_X1 U2416 ( .A(n3363), .ZN(n9019) );
  AOI22_X1 U2417 ( .A1(reg_mem[906]), .A2(n3361), .B1(n9025), .B2(data_w[2]), 
        .ZN(n3363) );
  INV_X1 U2418 ( .A(n3364), .ZN(n9020) );
  AOI22_X1 U2419 ( .A1(reg_mem[907]), .A2(n3361), .B1(n9025), .B2(data_w[3]), 
        .ZN(n3364) );
  INV_X1 U2420 ( .A(n3365), .ZN(n9021) );
  AOI22_X1 U2421 ( .A1(reg_mem[908]), .A2(n3361), .B1(n9025), .B2(data_w[4]), 
        .ZN(n3365) );
  INV_X1 U2422 ( .A(n3366), .ZN(n9022) );
  AOI22_X1 U2423 ( .A1(reg_mem[909]), .A2(n3361), .B1(n9025), .B2(data_w[5]), 
        .ZN(n3366) );
  INV_X1 U2424 ( .A(n3367), .ZN(n9023) );
  AOI22_X1 U2425 ( .A1(reg_mem[910]), .A2(n3361), .B1(n9025), .B2(data_w[6]), 
        .ZN(n3367) );
  INV_X1 U2426 ( .A(n3368), .ZN(n9024) );
  AOI22_X1 U2427 ( .A1(reg_mem[911]), .A2(n3361), .B1(n9025), .B2(data_w[7]), 
        .ZN(n3368) );
  INV_X1 U2428 ( .A(n3369), .ZN(n7864) );
  AOI22_X1 U2429 ( .A1(reg_mem[912]), .A2(n3370), .B1(n7872), .B2(data_w[0]), 
        .ZN(n3369) );
  INV_X1 U2430 ( .A(n3371), .ZN(n7865) );
  AOI22_X1 U2431 ( .A1(reg_mem[913]), .A2(n3370), .B1(n7872), .B2(data_w[1]), 
        .ZN(n3371) );
  INV_X1 U2432 ( .A(n3372), .ZN(n7866) );
  AOI22_X1 U2433 ( .A1(reg_mem[914]), .A2(n3370), .B1(n7872), .B2(data_w[2]), 
        .ZN(n3372) );
  INV_X1 U2434 ( .A(n3373), .ZN(n7867) );
  AOI22_X1 U2435 ( .A1(reg_mem[915]), .A2(n3370), .B1(n7872), .B2(data_w[3]), 
        .ZN(n3373) );
  INV_X1 U2436 ( .A(n3374), .ZN(n7868) );
  AOI22_X1 U2437 ( .A1(reg_mem[916]), .A2(n3370), .B1(n7872), .B2(data_w[4]), 
        .ZN(n3374) );
  INV_X1 U2438 ( .A(n3375), .ZN(n7869) );
  AOI22_X1 U2439 ( .A1(reg_mem[917]), .A2(n3370), .B1(n7872), .B2(data_w[5]), 
        .ZN(n3375) );
  INV_X1 U2440 ( .A(n3376), .ZN(n7870) );
  AOI22_X1 U2441 ( .A1(reg_mem[918]), .A2(n3370), .B1(n7872), .B2(data_w[6]), 
        .ZN(n3376) );
  INV_X1 U2442 ( .A(n3377), .ZN(n7871) );
  AOI22_X1 U2443 ( .A1(reg_mem[919]), .A2(n3370), .B1(n7872), .B2(data_w[7]), 
        .ZN(n3377) );
  INV_X1 U2444 ( .A(n3378), .ZN(n8441) );
  AOI22_X1 U2445 ( .A1(reg_mem[920]), .A2(n3379), .B1(n8449), .B2(data_w[0]), 
        .ZN(n3378) );
  INV_X1 U2446 ( .A(n3380), .ZN(n8442) );
  AOI22_X1 U2447 ( .A1(reg_mem[921]), .A2(n3379), .B1(n8449), .B2(data_w[1]), 
        .ZN(n3380) );
  INV_X1 U2448 ( .A(n3381), .ZN(n8443) );
  AOI22_X1 U2449 ( .A1(reg_mem[922]), .A2(n3379), .B1(n8449), .B2(data_w[2]), 
        .ZN(n3381) );
  INV_X1 U2450 ( .A(n3382), .ZN(n8444) );
  AOI22_X1 U2451 ( .A1(reg_mem[923]), .A2(n3379), .B1(n8449), .B2(data_w[3]), 
        .ZN(n3382) );
  INV_X1 U2452 ( .A(n3383), .ZN(n8445) );
  AOI22_X1 U2453 ( .A1(reg_mem[924]), .A2(n3379), .B1(n8449), .B2(data_w[4]), 
        .ZN(n3383) );
  INV_X1 U2454 ( .A(n3384), .ZN(n8446) );
  AOI22_X1 U2455 ( .A1(reg_mem[925]), .A2(n3379), .B1(n8449), .B2(data_w[5]), 
        .ZN(n3384) );
  INV_X1 U2456 ( .A(n3385), .ZN(n8447) );
  AOI22_X1 U2457 ( .A1(reg_mem[926]), .A2(n3379), .B1(n8449), .B2(data_w[6]), 
        .ZN(n3385) );
  INV_X1 U2458 ( .A(n3386), .ZN(n8448) );
  AOI22_X1 U2459 ( .A1(reg_mem[927]), .A2(n3379), .B1(n8449), .B2(data_w[7]), 
        .ZN(n3386) );
  INV_X1 U2460 ( .A(n3387), .ZN(n7144) );
  AOI22_X1 U2461 ( .A1(reg_mem[928]), .A2(n3388), .B1(n7152), .B2(data_w[0]), 
        .ZN(n3387) );
  INV_X1 U2462 ( .A(n3389), .ZN(n7145) );
  AOI22_X1 U2463 ( .A1(reg_mem[929]), .A2(n3388), .B1(n7152), .B2(data_w[1]), 
        .ZN(n3389) );
  INV_X1 U2464 ( .A(n3390), .ZN(n7146) );
  AOI22_X1 U2465 ( .A1(reg_mem[930]), .A2(n3388), .B1(n7152), .B2(data_w[2]), 
        .ZN(n3390) );
  INV_X1 U2466 ( .A(n3391), .ZN(n7147) );
  AOI22_X1 U2467 ( .A1(reg_mem[931]), .A2(n3388), .B1(n7152), .B2(data_w[3]), 
        .ZN(n3391) );
  INV_X1 U2468 ( .A(n3392), .ZN(n7148) );
  AOI22_X1 U2469 ( .A1(reg_mem[932]), .A2(n3388), .B1(n7152), .B2(data_w[4]), 
        .ZN(n3392) );
  INV_X1 U2470 ( .A(n3393), .ZN(n7149) );
  AOI22_X1 U2471 ( .A1(reg_mem[933]), .A2(n3388), .B1(n7152), .B2(data_w[5]), 
        .ZN(n3393) );
  INV_X1 U2472 ( .A(n3394), .ZN(n7150) );
  AOI22_X1 U2473 ( .A1(reg_mem[934]), .A2(n3388), .B1(n7152), .B2(data_w[6]), 
        .ZN(n3394) );
  INV_X1 U2474 ( .A(n3395), .ZN(n7151) );
  AOI22_X1 U2475 ( .A1(reg_mem[935]), .A2(n3388), .B1(n7152), .B2(data_w[7]), 
        .ZN(n3395) );
  INV_X1 U2476 ( .A(n3396), .ZN(n8873) );
  AOI22_X1 U2477 ( .A1(reg_mem[936]), .A2(n3397), .B1(n8881), .B2(data_w[0]), 
        .ZN(n3396) );
  INV_X1 U2478 ( .A(n3398), .ZN(n8874) );
  AOI22_X1 U2479 ( .A1(reg_mem[937]), .A2(n3397), .B1(n8881), .B2(data_w[1]), 
        .ZN(n3398) );
  INV_X1 U2480 ( .A(n3399), .ZN(n8875) );
  AOI22_X1 U2481 ( .A1(reg_mem[938]), .A2(n3397), .B1(n8881), .B2(data_w[2]), 
        .ZN(n3399) );
  INV_X1 U2482 ( .A(n3400), .ZN(n8876) );
  AOI22_X1 U2483 ( .A1(reg_mem[939]), .A2(n3397), .B1(n8881), .B2(data_w[3]), 
        .ZN(n3400) );
  INV_X1 U2484 ( .A(n3401), .ZN(n8877) );
  AOI22_X1 U2485 ( .A1(reg_mem[940]), .A2(n3397), .B1(n8881), .B2(data_w[4]), 
        .ZN(n3401) );
  INV_X1 U2486 ( .A(n3402), .ZN(n8878) );
  AOI22_X1 U2487 ( .A1(reg_mem[941]), .A2(n3397), .B1(n8881), .B2(data_w[5]), 
        .ZN(n3402) );
  INV_X1 U2488 ( .A(n3403), .ZN(n8879) );
  AOI22_X1 U2489 ( .A1(reg_mem[942]), .A2(n3397), .B1(n8881), .B2(data_w[6]), 
        .ZN(n3403) );
  INV_X1 U2490 ( .A(n3404), .ZN(n8880) );
  AOI22_X1 U2491 ( .A1(reg_mem[943]), .A2(n3397), .B1(n8881), .B2(data_w[7]), 
        .ZN(n3404) );
  INV_X1 U2492 ( .A(n3405), .ZN(n7720) );
  AOI22_X1 U2493 ( .A1(reg_mem[944]), .A2(n3406), .B1(n7728), .B2(data_w[0]), 
        .ZN(n3405) );
  INV_X1 U2494 ( .A(n3407), .ZN(n7721) );
  AOI22_X1 U2495 ( .A1(reg_mem[945]), .A2(n3406), .B1(n7728), .B2(data_w[1]), 
        .ZN(n3407) );
  INV_X1 U2496 ( .A(n3408), .ZN(n7722) );
  AOI22_X1 U2497 ( .A1(reg_mem[946]), .A2(n3406), .B1(n7728), .B2(data_w[2]), 
        .ZN(n3408) );
  INV_X1 U2498 ( .A(n3409), .ZN(n7723) );
  AOI22_X1 U2499 ( .A1(reg_mem[947]), .A2(n3406), .B1(n7728), .B2(data_w[3]), 
        .ZN(n3409) );
  INV_X1 U2500 ( .A(n3410), .ZN(n7724) );
  AOI22_X1 U2501 ( .A1(reg_mem[948]), .A2(n3406), .B1(n7728), .B2(data_w[4]), 
        .ZN(n3410) );
  INV_X1 U2502 ( .A(n3411), .ZN(n7725) );
  AOI22_X1 U2503 ( .A1(reg_mem[949]), .A2(n3406), .B1(n7728), .B2(data_w[5]), 
        .ZN(n3411) );
  INV_X1 U2504 ( .A(n3412), .ZN(n7726) );
  AOI22_X1 U2505 ( .A1(reg_mem[950]), .A2(n3406), .B1(n7728), .B2(data_w[6]), 
        .ZN(n3412) );
  INV_X1 U2506 ( .A(n3413), .ZN(n7727) );
  AOI22_X1 U2507 ( .A1(reg_mem[951]), .A2(n3406), .B1(n7728), .B2(data_w[7]), 
        .ZN(n3413) );
  INV_X1 U2508 ( .A(n3414), .ZN(n8297) );
  AOI22_X1 U2509 ( .A1(reg_mem[952]), .A2(n3415), .B1(n8305), .B2(data_w[0]), 
        .ZN(n3414) );
  INV_X1 U2510 ( .A(n3416), .ZN(n8298) );
  AOI22_X1 U2511 ( .A1(reg_mem[953]), .A2(n3415), .B1(n8305), .B2(data_w[1]), 
        .ZN(n3416) );
  INV_X1 U2512 ( .A(n3417), .ZN(n8299) );
  AOI22_X1 U2513 ( .A1(reg_mem[954]), .A2(n3415), .B1(n8305), .B2(data_w[2]), 
        .ZN(n3417) );
  INV_X1 U2514 ( .A(n3418), .ZN(n8300) );
  AOI22_X1 U2515 ( .A1(reg_mem[955]), .A2(n3415), .B1(n8305), .B2(data_w[3]), 
        .ZN(n3418) );
  INV_X1 U2516 ( .A(n3419), .ZN(n8301) );
  AOI22_X1 U2517 ( .A1(reg_mem[956]), .A2(n3415), .B1(n8305), .B2(data_w[4]), 
        .ZN(n3419) );
  INV_X1 U2518 ( .A(n3420), .ZN(n8302) );
  AOI22_X1 U2519 ( .A1(reg_mem[957]), .A2(n3415), .B1(n8305), .B2(data_w[5]), 
        .ZN(n3420) );
  INV_X1 U2520 ( .A(n3421), .ZN(n8303) );
  AOI22_X1 U2521 ( .A1(reg_mem[958]), .A2(n3415), .B1(n8305), .B2(data_w[6]), 
        .ZN(n3421) );
  INV_X1 U2522 ( .A(n3422), .ZN(n8304) );
  AOI22_X1 U2523 ( .A1(reg_mem[959]), .A2(n3415), .B1(n8305), .B2(data_w[7]), 
        .ZN(n3422) );
  INV_X1 U2524 ( .A(n3423), .ZN(n7000) );
  AOI22_X1 U2525 ( .A1(reg_mem[960]), .A2(n3424), .B1(n7008), .B2(data_w[0]), 
        .ZN(n3423) );
  INV_X1 U2526 ( .A(n3425), .ZN(n7001) );
  AOI22_X1 U2527 ( .A1(reg_mem[961]), .A2(n3424), .B1(n7008), .B2(data_w[1]), 
        .ZN(n3425) );
  INV_X1 U2528 ( .A(n3426), .ZN(n7002) );
  AOI22_X1 U2529 ( .A1(reg_mem[962]), .A2(n3424), .B1(n7008), .B2(data_w[2]), 
        .ZN(n3426) );
  INV_X1 U2530 ( .A(n3427), .ZN(n7003) );
  AOI22_X1 U2531 ( .A1(reg_mem[963]), .A2(n3424), .B1(n7008), .B2(data_w[3]), 
        .ZN(n3427) );
  INV_X1 U2532 ( .A(n3428), .ZN(n7004) );
  AOI22_X1 U2533 ( .A1(reg_mem[964]), .A2(n3424), .B1(n7008), .B2(data_w[4]), 
        .ZN(n3428) );
  INV_X1 U2534 ( .A(n3429), .ZN(n7005) );
  AOI22_X1 U2535 ( .A1(reg_mem[965]), .A2(n3424), .B1(n7008), .B2(data_w[5]), 
        .ZN(n3429) );
  INV_X1 U2536 ( .A(n3430), .ZN(n7006) );
  AOI22_X1 U2537 ( .A1(reg_mem[966]), .A2(n3424), .B1(n7008), .B2(data_w[6]), 
        .ZN(n3430) );
  INV_X1 U2538 ( .A(n3431), .ZN(n7007) );
  AOI22_X1 U2539 ( .A1(reg_mem[967]), .A2(n3424), .B1(n7008), .B2(data_w[7]), 
        .ZN(n3431) );
  INV_X1 U2540 ( .A(n3432), .ZN(n8729) );
  AOI22_X1 U2541 ( .A1(reg_mem[968]), .A2(n3433), .B1(n8737), .B2(data_w[0]), 
        .ZN(n3432) );
  INV_X1 U2542 ( .A(n3434), .ZN(n8730) );
  AOI22_X1 U2543 ( .A1(reg_mem[969]), .A2(n3433), .B1(n8737), .B2(data_w[1]), 
        .ZN(n3434) );
  INV_X1 U2544 ( .A(n3435), .ZN(n8731) );
  AOI22_X1 U2545 ( .A1(reg_mem[970]), .A2(n3433), .B1(n8737), .B2(data_w[2]), 
        .ZN(n3435) );
  INV_X1 U2546 ( .A(n3436), .ZN(n8732) );
  AOI22_X1 U2547 ( .A1(reg_mem[971]), .A2(n3433), .B1(n8737), .B2(data_w[3]), 
        .ZN(n3436) );
  INV_X1 U2548 ( .A(n3437), .ZN(n8733) );
  AOI22_X1 U2549 ( .A1(reg_mem[972]), .A2(n3433), .B1(n8737), .B2(data_w[4]), 
        .ZN(n3437) );
  INV_X1 U2550 ( .A(n3438), .ZN(n8734) );
  AOI22_X1 U2551 ( .A1(reg_mem[973]), .A2(n3433), .B1(n8737), .B2(data_w[5]), 
        .ZN(n3438) );
  INV_X1 U2552 ( .A(n3439), .ZN(n8735) );
  AOI22_X1 U2553 ( .A1(reg_mem[974]), .A2(n3433), .B1(n8737), .B2(data_w[6]), 
        .ZN(n3439) );
  INV_X1 U2554 ( .A(n3440), .ZN(n8736) );
  AOI22_X1 U2555 ( .A1(reg_mem[975]), .A2(n3433), .B1(n8737), .B2(data_w[7]), 
        .ZN(n3440) );
  INV_X1 U2556 ( .A(n3441), .ZN(n7576) );
  AOI22_X1 U2557 ( .A1(reg_mem[976]), .A2(n3442), .B1(n7584), .B2(data_w[0]), 
        .ZN(n3441) );
  INV_X1 U2558 ( .A(n3443), .ZN(n7577) );
  AOI22_X1 U2559 ( .A1(reg_mem[977]), .A2(n3442), .B1(n7584), .B2(data_w[1]), 
        .ZN(n3443) );
  INV_X1 U2560 ( .A(n3444), .ZN(n7578) );
  AOI22_X1 U2561 ( .A1(reg_mem[978]), .A2(n3442), .B1(n7584), .B2(data_w[2]), 
        .ZN(n3444) );
  INV_X1 U2562 ( .A(n3445), .ZN(n7579) );
  AOI22_X1 U2563 ( .A1(reg_mem[979]), .A2(n3442), .B1(n7584), .B2(data_w[3]), 
        .ZN(n3445) );
  INV_X1 U2564 ( .A(n3446), .ZN(n7580) );
  AOI22_X1 U2565 ( .A1(reg_mem[980]), .A2(n3442), .B1(n7584), .B2(data_w[4]), 
        .ZN(n3446) );
  INV_X1 U2566 ( .A(n3447), .ZN(n7581) );
  AOI22_X1 U2567 ( .A1(reg_mem[981]), .A2(n3442), .B1(n7584), .B2(data_w[5]), 
        .ZN(n3447) );
  INV_X1 U2568 ( .A(n3448), .ZN(n7582) );
  AOI22_X1 U2569 ( .A1(reg_mem[982]), .A2(n3442), .B1(n7584), .B2(data_w[6]), 
        .ZN(n3448) );
  INV_X1 U2570 ( .A(n3449), .ZN(n7583) );
  AOI22_X1 U2571 ( .A1(reg_mem[983]), .A2(n3442), .B1(n7584), .B2(data_w[7]), 
        .ZN(n3449) );
  INV_X1 U2572 ( .A(n3450), .ZN(n8153) );
  AOI22_X1 U2573 ( .A1(reg_mem[984]), .A2(n3451), .B1(n8161), .B2(data_w[0]), 
        .ZN(n3450) );
  INV_X1 U2574 ( .A(n3452), .ZN(n8154) );
  AOI22_X1 U2575 ( .A1(reg_mem[985]), .A2(n3451), .B1(n8161), .B2(data_w[1]), 
        .ZN(n3452) );
  INV_X1 U2576 ( .A(n3453), .ZN(n8155) );
  AOI22_X1 U2577 ( .A1(reg_mem[986]), .A2(n3451), .B1(n8161), .B2(data_w[2]), 
        .ZN(n3453) );
  INV_X1 U2578 ( .A(n3454), .ZN(n8156) );
  AOI22_X1 U2579 ( .A1(reg_mem[987]), .A2(n3451), .B1(n8161), .B2(data_w[3]), 
        .ZN(n3454) );
  INV_X1 U2580 ( .A(n3455), .ZN(n8157) );
  AOI22_X1 U2581 ( .A1(reg_mem[988]), .A2(n3451), .B1(n8161), .B2(data_w[4]), 
        .ZN(n3455) );
  INV_X1 U2582 ( .A(n3456), .ZN(n8158) );
  AOI22_X1 U2583 ( .A1(reg_mem[989]), .A2(n3451), .B1(n8161), .B2(data_w[5]), 
        .ZN(n3456) );
  INV_X1 U2584 ( .A(n3457), .ZN(n8159) );
  AOI22_X1 U2585 ( .A1(reg_mem[990]), .A2(n3451), .B1(n8161), .B2(data_w[6]), 
        .ZN(n3457) );
  INV_X1 U2586 ( .A(n3458), .ZN(n8160) );
  AOI22_X1 U2587 ( .A1(reg_mem[991]), .A2(n3451), .B1(n8161), .B2(data_w[7]), 
        .ZN(n3458) );
  INV_X1 U2588 ( .A(n3895), .ZN(n6829) );
  AOI22_X1 U2589 ( .A1(reg_mem[1376]), .A2(n3896), .B1(n6837), .B2(data_w[0]), 
        .ZN(n3895) );
  INV_X1 U2590 ( .A(n3897), .ZN(n6830) );
  AOI22_X1 U2591 ( .A1(reg_mem[1377]), .A2(n3896), .B1(n6837), .B2(data_w[1]), 
        .ZN(n3897) );
  INV_X1 U2592 ( .A(n3898), .ZN(n6831) );
  AOI22_X1 U2593 ( .A1(reg_mem[1378]), .A2(n3896), .B1(n6837), .B2(data_w[2]), 
        .ZN(n3898) );
  INV_X1 U2594 ( .A(n3899), .ZN(n6832) );
  AOI22_X1 U2595 ( .A1(reg_mem[1379]), .A2(n3896), .B1(n6837), .B2(data_w[3]), 
        .ZN(n3899) );
  INV_X1 U2596 ( .A(n3900), .ZN(n6833) );
  AOI22_X1 U2597 ( .A1(reg_mem[1380]), .A2(n3896), .B1(n6837), .B2(data_w[4]), 
        .ZN(n3900) );
  INV_X1 U2598 ( .A(n3901), .ZN(n6834) );
  AOI22_X1 U2599 ( .A1(reg_mem[1381]), .A2(n3896), .B1(n6837), .B2(data_w[5]), 
        .ZN(n3901) );
  INV_X1 U2600 ( .A(n3902), .ZN(n6835) );
  AOI22_X1 U2601 ( .A1(reg_mem[1382]), .A2(n3896), .B1(n6837), .B2(data_w[6]), 
        .ZN(n3902) );
  INV_X1 U2602 ( .A(n3903), .ZN(n6836) );
  AOI22_X1 U2603 ( .A1(reg_mem[1383]), .A2(n3896), .B1(n6837), .B2(data_w[7]), 
        .ZN(n3903) );
  INV_X1 U2604 ( .A(n3904), .ZN(n8558) );
  AOI22_X1 U2605 ( .A1(reg_mem[1384]), .A2(n3905), .B1(n8566), .B2(data_w[0]), 
        .ZN(n3904) );
  INV_X1 U2606 ( .A(n3906), .ZN(n8559) );
  AOI22_X1 U2607 ( .A1(reg_mem[1385]), .A2(n3905), .B1(n8566), .B2(data_w[1]), 
        .ZN(n3906) );
  INV_X1 U2608 ( .A(n3907), .ZN(n8560) );
  AOI22_X1 U2609 ( .A1(reg_mem[1386]), .A2(n3905), .B1(n8566), .B2(data_w[2]), 
        .ZN(n3907) );
  INV_X1 U2610 ( .A(n3908), .ZN(n8561) );
  AOI22_X1 U2611 ( .A1(reg_mem[1387]), .A2(n3905), .B1(n8566), .B2(data_w[3]), 
        .ZN(n3908) );
  INV_X1 U2612 ( .A(n3909), .ZN(n8562) );
  AOI22_X1 U2613 ( .A1(reg_mem[1388]), .A2(n3905), .B1(n8566), .B2(data_w[4]), 
        .ZN(n3909) );
  INV_X1 U2614 ( .A(n3910), .ZN(n8563) );
  AOI22_X1 U2615 ( .A1(reg_mem[1389]), .A2(n3905), .B1(n8566), .B2(data_w[5]), 
        .ZN(n3910) );
  INV_X1 U2616 ( .A(n3911), .ZN(n8564) );
  AOI22_X1 U2617 ( .A1(reg_mem[1390]), .A2(n3905), .B1(n8566), .B2(data_w[6]), 
        .ZN(n3911) );
  INV_X1 U2618 ( .A(n3912), .ZN(n8565) );
  AOI22_X1 U2619 ( .A1(reg_mem[1391]), .A2(n3905), .B1(n8566), .B2(data_w[7]), 
        .ZN(n3912) );
  INV_X1 U2620 ( .A(n3913), .ZN(n7405) );
  AOI22_X1 U2621 ( .A1(reg_mem[1392]), .A2(n3914), .B1(n7413), .B2(data_w[0]), 
        .ZN(n3913) );
  INV_X1 U2622 ( .A(n3915), .ZN(n7406) );
  AOI22_X1 U2623 ( .A1(reg_mem[1393]), .A2(n3914), .B1(n7413), .B2(data_w[1]), 
        .ZN(n3915) );
  INV_X1 U2624 ( .A(n3916), .ZN(n7407) );
  AOI22_X1 U2625 ( .A1(reg_mem[1394]), .A2(n3914), .B1(n7413), .B2(data_w[2]), 
        .ZN(n3916) );
  INV_X1 U2626 ( .A(n3917), .ZN(n7408) );
  AOI22_X1 U2627 ( .A1(reg_mem[1395]), .A2(n3914), .B1(n7413), .B2(data_w[3]), 
        .ZN(n3917) );
  INV_X1 U2628 ( .A(n3918), .ZN(n7409) );
  AOI22_X1 U2629 ( .A1(reg_mem[1396]), .A2(n3914), .B1(n7413), .B2(data_w[4]), 
        .ZN(n3918) );
  INV_X1 U2630 ( .A(n3919), .ZN(n7410) );
  AOI22_X1 U2631 ( .A1(reg_mem[1397]), .A2(n3914), .B1(n7413), .B2(data_w[5]), 
        .ZN(n3919) );
  INV_X1 U2632 ( .A(n3920), .ZN(n7411) );
  AOI22_X1 U2633 ( .A1(reg_mem[1398]), .A2(n3914), .B1(n7413), .B2(data_w[6]), 
        .ZN(n3920) );
  INV_X1 U2634 ( .A(n3921), .ZN(n7412) );
  AOI22_X1 U2635 ( .A1(reg_mem[1399]), .A2(n3914), .B1(n7413), .B2(data_w[7]), 
        .ZN(n3921) );
  INV_X1 U2636 ( .A(n3922), .ZN(n7982) );
  AOI22_X1 U2637 ( .A1(reg_mem[1400]), .A2(n3923), .B1(n7990), .B2(data_w[0]), 
        .ZN(n3922) );
  INV_X1 U2638 ( .A(n3924), .ZN(n7983) );
  AOI22_X1 U2639 ( .A1(reg_mem[1401]), .A2(n3923), .B1(n7990), .B2(data_w[1]), 
        .ZN(n3924) );
  INV_X1 U2640 ( .A(n3925), .ZN(n7984) );
  AOI22_X1 U2641 ( .A1(reg_mem[1402]), .A2(n3923), .B1(n7990), .B2(data_w[2]), 
        .ZN(n3925) );
  INV_X1 U2642 ( .A(n3926), .ZN(n7985) );
  AOI22_X1 U2643 ( .A1(reg_mem[1403]), .A2(n3923), .B1(n7990), .B2(data_w[3]), 
        .ZN(n3926) );
  INV_X1 U2644 ( .A(n3927), .ZN(n7986) );
  AOI22_X1 U2645 ( .A1(reg_mem[1404]), .A2(n3923), .B1(n7990), .B2(data_w[4]), 
        .ZN(n3927) );
  INV_X1 U2646 ( .A(n3928), .ZN(n7987) );
  AOI22_X1 U2647 ( .A1(reg_mem[1405]), .A2(n3923), .B1(n7990), .B2(data_w[5]), 
        .ZN(n3928) );
  INV_X1 U2648 ( .A(n3929), .ZN(n7988) );
  AOI22_X1 U2649 ( .A1(reg_mem[1406]), .A2(n3923), .B1(n7990), .B2(data_w[6]), 
        .ZN(n3929) );
  INV_X1 U2650 ( .A(n3930), .ZN(n7989) );
  AOI22_X1 U2651 ( .A1(reg_mem[1407]), .A2(n3923), .B1(n7990), .B2(data_w[7]), 
        .ZN(n3930) );
  INV_X1 U2652 ( .A(n3931), .ZN(n7252) );
  AOI22_X1 U2653 ( .A1(reg_mem[1408]), .A2(n3932), .B1(n7260), .B2(data_w[0]), 
        .ZN(n3931) );
  INV_X1 U2654 ( .A(n3933), .ZN(n7253) );
  AOI22_X1 U2655 ( .A1(reg_mem[1409]), .A2(n3932), .B1(n7260), .B2(data_w[1]), 
        .ZN(n3933) );
  INV_X1 U2656 ( .A(n3934), .ZN(n7254) );
  AOI22_X1 U2657 ( .A1(reg_mem[1410]), .A2(n3932), .B1(n7260), .B2(data_w[2]), 
        .ZN(n3934) );
  INV_X1 U2658 ( .A(n3935), .ZN(n7255) );
  AOI22_X1 U2659 ( .A1(reg_mem[1411]), .A2(n3932), .B1(n7260), .B2(data_w[3]), 
        .ZN(n3935) );
  INV_X1 U2660 ( .A(n3936), .ZN(n7256) );
  AOI22_X1 U2661 ( .A1(reg_mem[1412]), .A2(n3932), .B1(n7260), .B2(data_w[4]), 
        .ZN(n3936) );
  INV_X1 U2662 ( .A(n3937), .ZN(n7257) );
  AOI22_X1 U2663 ( .A1(reg_mem[1413]), .A2(n3932), .B1(n7260), .B2(data_w[5]), 
        .ZN(n3937) );
  INV_X1 U2664 ( .A(n3938), .ZN(n7258) );
  AOI22_X1 U2665 ( .A1(reg_mem[1414]), .A2(n3932), .B1(n7260), .B2(data_w[6]), 
        .ZN(n3938) );
  INV_X1 U2666 ( .A(n3939), .ZN(n7259) );
  AOI22_X1 U2667 ( .A1(reg_mem[1415]), .A2(n3932), .B1(n7260), .B2(data_w[7]), 
        .ZN(n3939) );
  INV_X1 U2668 ( .A(n3941), .ZN(n8981) );
  AOI22_X1 U2669 ( .A1(reg_mem[1416]), .A2(n3942), .B1(n8989), .B2(data_w[0]), 
        .ZN(n3941) );
  INV_X1 U2670 ( .A(n3943), .ZN(n8982) );
  AOI22_X1 U2671 ( .A1(reg_mem[1417]), .A2(n3942), .B1(n8989), .B2(data_w[1]), 
        .ZN(n3943) );
  INV_X1 U2672 ( .A(n3944), .ZN(n8983) );
  AOI22_X1 U2673 ( .A1(reg_mem[1418]), .A2(n3942), .B1(n8989), .B2(data_w[2]), 
        .ZN(n3944) );
  INV_X1 U2674 ( .A(n3945), .ZN(n8984) );
  AOI22_X1 U2675 ( .A1(reg_mem[1419]), .A2(n3942), .B1(n8989), .B2(data_w[3]), 
        .ZN(n3945) );
  INV_X1 U2676 ( .A(n3946), .ZN(n8985) );
  AOI22_X1 U2677 ( .A1(reg_mem[1420]), .A2(n3942), .B1(n8989), .B2(data_w[4]), 
        .ZN(n3946) );
  INV_X1 U2678 ( .A(n3947), .ZN(n8986) );
  AOI22_X1 U2679 ( .A1(reg_mem[1421]), .A2(n3942), .B1(n8989), .B2(data_w[5]), 
        .ZN(n3947) );
  INV_X1 U2680 ( .A(n3948), .ZN(n8987) );
  AOI22_X1 U2681 ( .A1(reg_mem[1422]), .A2(n3942), .B1(n8989), .B2(data_w[6]), 
        .ZN(n3948) );
  INV_X1 U2682 ( .A(n3949), .ZN(n8988) );
  AOI22_X1 U2683 ( .A1(reg_mem[1423]), .A2(n3942), .B1(n8989), .B2(data_w[7]), 
        .ZN(n3949) );
  INV_X1 U2684 ( .A(n3950), .ZN(n7828) );
  AOI22_X1 U2685 ( .A1(reg_mem[1424]), .A2(n3951), .B1(n7836), .B2(data_w[0]), 
        .ZN(n3950) );
  INV_X1 U2686 ( .A(n3952), .ZN(n7829) );
  AOI22_X1 U2687 ( .A1(reg_mem[1425]), .A2(n3951), .B1(n7836), .B2(data_w[1]), 
        .ZN(n3952) );
  INV_X1 U2688 ( .A(n3953), .ZN(n7830) );
  AOI22_X1 U2689 ( .A1(reg_mem[1426]), .A2(n3951), .B1(n7836), .B2(data_w[2]), 
        .ZN(n3953) );
  INV_X1 U2690 ( .A(n3954), .ZN(n7831) );
  AOI22_X1 U2691 ( .A1(reg_mem[1427]), .A2(n3951), .B1(n7836), .B2(data_w[3]), 
        .ZN(n3954) );
  INV_X1 U2692 ( .A(n3955), .ZN(n7832) );
  AOI22_X1 U2693 ( .A1(reg_mem[1428]), .A2(n3951), .B1(n7836), .B2(data_w[4]), 
        .ZN(n3955) );
  INV_X1 U2694 ( .A(n3956), .ZN(n7833) );
  AOI22_X1 U2695 ( .A1(reg_mem[1429]), .A2(n3951), .B1(n7836), .B2(data_w[5]), 
        .ZN(n3956) );
  INV_X1 U2696 ( .A(n3957), .ZN(n7834) );
  AOI22_X1 U2697 ( .A1(reg_mem[1430]), .A2(n3951), .B1(n7836), .B2(data_w[6]), 
        .ZN(n3957) );
  INV_X1 U2698 ( .A(n3958), .ZN(n7835) );
  AOI22_X1 U2699 ( .A1(reg_mem[1431]), .A2(n3951), .B1(n7836), .B2(data_w[7]), 
        .ZN(n3958) );
  INV_X1 U2700 ( .A(n3959), .ZN(n8405) );
  AOI22_X1 U2701 ( .A1(reg_mem[1432]), .A2(n3960), .B1(n8413), .B2(data_w[0]), 
        .ZN(n3959) );
  INV_X1 U2702 ( .A(n3961), .ZN(n8406) );
  AOI22_X1 U2703 ( .A1(reg_mem[1433]), .A2(n3960), .B1(n8413), .B2(data_w[1]), 
        .ZN(n3961) );
  INV_X1 U2704 ( .A(n3962), .ZN(n8407) );
  AOI22_X1 U2705 ( .A1(reg_mem[1434]), .A2(n3960), .B1(n8413), .B2(data_w[2]), 
        .ZN(n3962) );
  INV_X1 U2706 ( .A(n3963), .ZN(n8408) );
  AOI22_X1 U2707 ( .A1(reg_mem[1435]), .A2(n3960), .B1(n8413), .B2(data_w[3]), 
        .ZN(n3963) );
  INV_X1 U2708 ( .A(n3964), .ZN(n8409) );
  AOI22_X1 U2709 ( .A1(reg_mem[1436]), .A2(n3960), .B1(n8413), .B2(data_w[4]), 
        .ZN(n3964) );
  INV_X1 U2710 ( .A(n3965), .ZN(n8410) );
  AOI22_X1 U2711 ( .A1(reg_mem[1437]), .A2(n3960), .B1(n8413), .B2(data_w[5]), 
        .ZN(n3965) );
  INV_X1 U2712 ( .A(n3966), .ZN(n8411) );
  AOI22_X1 U2713 ( .A1(reg_mem[1438]), .A2(n3960), .B1(n8413), .B2(data_w[6]), 
        .ZN(n3966) );
  INV_X1 U2714 ( .A(n3967), .ZN(n8412) );
  AOI22_X1 U2715 ( .A1(reg_mem[1439]), .A2(n3960), .B1(n8413), .B2(data_w[7]), 
        .ZN(n3967) );
  INV_X1 U2716 ( .A(n3968), .ZN(n7108) );
  AOI22_X1 U2717 ( .A1(reg_mem[1440]), .A2(n3969), .B1(n7116), .B2(data_w[0]), 
        .ZN(n3968) );
  INV_X1 U2718 ( .A(n3970), .ZN(n7109) );
  AOI22_X1 U2719 ( .A1(reg_mem[1441]), .A2(n3969), .B1(n7116), .B2(data_w[1]), 
        .ZN(n3970) );
  INV_X1 U2720 ( .A(n3971), .ZN(n7110) );
  AOI22_X1 U2721 ( .A1(reg_mem[1442]), .A2(n3969), .B1(n7116), .B2(data_w[2]), 
        .ZN(n3971) );
  INV_X1 U2722 ( .A(n3972), .ZN(n7111) );
  AOI22_X1 U2723 ( .A1(reg_mem[1443]), .A2(n3969), .B1(n7116), .B2(data_w[3]), 
        .ZN(n3972) );
  INV_X1 U2724 ( .A(n3973), .ZN(n7112) );
  AOI22_X1 U2725 ( .A1(reg_mem[1444]), .A2(n3969), .B1(n7116), .B2(data_w[4]), 
        .ZN(n3973) );
  INV_X1 U2726 ( .A(n3974), .ZN(n7113) );
  AOI22_X1 U2727 ( .A1(reg_mem[1445]), .A2(n3969), .B1(n7116), .B2(data_w[5]), 
        .ZN(n3974) );
  INV_X1 U2728 ( .A(n3975), .ZN(n7114) );
  AOI22_X1 U2729 ( .A1(reg_mem[1446]), .A2(n3969), .B1(n7116), .B2(data_w[6]), 
        .ZN(n3975) );
  INV_X1 U2730 ( .A(n3976), .ZN(n7115) );
  AOI22_X1 U2731 ( .A1(reg_mem[1447]), .A2(n3969), .B1(n7116), .B2(data_w[7]), 
        .ZN(n3976) );
  INV_X1 U2732 ( .A(n3977), .ZN(n8837) );
  AOI22_X1 U2733 ( .A1(reg_mem[1448]), .A2(n3978), .B1(n8845), .B2(data_w[0]), 
        .ZN(n3977) );
  INV_X1 U2734 ( .A(n3979), .ZN(n8838) );
  AOI22_X1 U2735 ( .A1(reg_mem[1449]), .A2(n3978), .B1(n8845), .B2(data_w[1]), 
        .ZN(n3979) );
  INV_X1 U2736 ( .A(n3980), .ZN(n8839) );
  AOI22_X1 U2737 ( .A1(reg_mem[1450]), .A2(n3978), .B1(n8845), .B2(data_w[2]), 
        .ZN(n3980) );
  INV_X1 U2738 ( .A(n3981), .ZN(n8840) );
  AOI22_X1 U2739 ( .A1(reg_mem[1451]), .A2(n3978), .B1(n8845), .B2(data_w[3]), 
        .ZN(n3981) );
  INV_X1 U2740 ( .A(n3982), .ZN(n8841) );
  AOI22_X1 U2741 ( .A1(reg_mem[1452]), .A2(n3978), .B1(n8845), .B2(data_w[4]), 
        .ZN(n3982) );
  INV_X1 U2742 ( .A(n3983), .ZN(n8842) );
  AOI22_X1 U2743 ( .A1(reg_mem[1453]), .A2(n3978), .B1(n8845), .B2(data_w[5]), 
        .ZN(n3983) );
  INV_X1 U2744 ( .A(n3984), .ZN(n8843) );
  AOI22_X1 U2745 ( .A1(reg_mem[1454]), .A2(n3978), .B1(n8845), .B2(data_w[6]), 
        .ZN(n3984) );
  INV_X1 U2746 ( .A(n3985), .ZN(n8844) );
  AOI22_X1 U2747 ( .A1(reg_mem[1455]), .A2(n3978), .B1(n8845), .B2(data_w[7]), 
        .ZN(n3985) );
  INV_X1 U2748 ( .A(n3986), .ZN(n7684) );
  AOI22_X1 U2749 ( .A1(reg_mem[1456]), .A2(n3987), .B1(n7692), .B2(data_w[0]), 
        .ZN(n3986) );
  INV_X1 U2750 ( .A(n3988), .ZN(n7685) );
  AOI22_X1 U2751 ( .A1(reg_mem[1457]), .A2(n3987), .B1(n7692), .B2(data_w[1]), 
        .ZN(n3988) );
  INV_X1 U2752 ( .A(n3989), .ZN(n7686) );
  AOI22_X1 U2753 ( .A1(reg_mem[1458]), .A2(n3987), .B1(n7692), .B2(data_w[2]), 
        .ZN(n3989) );
  INV_X1 U2754 ( .A(n3990), .ZN(n7687) );
  AOI22_X1 U2755 ( .A1(reg_mem[1459]), .A2(n3987), .B1(n7692), .B2(data_w[3]), 
        .ZN(n3990) );
  INV_X1 U2756 ( .A(n3991), .ZN(n7688) );
  AOI22_X1 U2757 ( .A1(reg_mem[1460]), .A2(n3987), .B1(n7692), .B2(data_w[4]), 
        .ZN(n3991) );
  INV_X1 U2758 ( .A(n3992), .ZN(n7689) );
  AOI22_X1 U2759 ( .A1(reg_mem[1461]), .A2(n3987), .B1(n7692), .B2(data_w[5]), 
        .ZN(n3992) );
  INV_X1 U2760 ( .A(n3993), .ZN(n7690) );
  AOI22_X1 U2761 ( .A1(reg_mem[1462]), .A2(n3987), .B1(n7692), .B2(data_w[6]), 
        .ZN(n3993) );
  INV_X1 U2762 ( .A(n3994), .ZN(n7691) );
  AOI22_X1 U2763 ( .A1(reg_mem[1463]), .A2(n3987), .B1(n7692), .B2(data_w[7]), 
        .ZN(n3994) );
  INV_X1 U2764 ( .A(n3995), .ZN(n8261) );
  AOI22_X1 U2765 ( .A1(reg_mem[1464]), .A2(n3996), .B1(n8269), .B2(data_w[0]), 
        .ZN(n3995) );
  INV_X1 U2766 ( .A(n3997), .ZN(n8262) );
  AOI22_X1 U2767 ( .A1(reg_mem[1465]), .A2(n3996), .B1(n8269), .B2(data_w[1]), 
        .ZN(n3997) );
  INV_X1 U2768 ( .A(n3998), .ZN(n8263) );
  AOI22_X1 U2769 ( .A1(reg_mem[1466]), .A2(n3996), .B1(n8269), .B2(data_w[2]), 
        .ZN(n3998) );
  INV_X1 U2770 ( .A(n3999), .ZN(n8264) );
  AOI22_X1 U2771 ( .A1(reg_mem[1467]), .A2(n3996), .B1(n8269), .B2(data_w[3]), 
        .ZN(n3999) );
  INV_X1 U2772 ( .A(n4000), .ZN(n8265) );
  AOI22_X1 U2773 ( .A1(reg_mem[1468]), .A2(n3996), .B1(n8269), .B2(data_w[4]), 
        .ZN(n4000) );
  INV_X1 U2774 ( .A(n4001), .ZN(n8266) );
  AOI22_X1 U2775 ( .A1(reg_mem[1469]), .A2(n3996), .B1(n8269), .B2(data_w[5]), 
        .ZN(n4001) );
  INV_X1 U2776 ( .A(n4002), .ZN(n8267) );
  AOI22_X1 U2777 ( .A1(reg_mem[1470]), .A2(n3996), .B1(n8269), .B2(data_w[6]), 
        .ZN(n4002) );
  INV_X1 U2778 ( .A(n4003), .ZN(n8268) );
  AOI22_X1 U2779 ( .A1(reg_mem[1471]), .A2(n3996), .B1(n8269), .B2(data_w[7]), 
        .ZN(n4003) );
  INV_X1 U2780 ( .A(n4004), .ZN(n6964) );
  AOI22_X1 U2781 ( .A1(reg_mem[1472]), .A2(n4005), .B1(n6972), .B2(data_w[0]), 
        .ZN(n4004) );
  INV_X1 U2782 ( .A(n4006), .ZN(n6965) );
  AOI22_X1 U2783 ( .A1(reg_mem[1473]), .A2(n4005), .B1(n6972), .B2(data_w[1]), 
        .ZN(n4006) );
  INV_X1 U2784 ( .A(n4007), .ZN(n6966) );
  AOI22_X1 U2785 ( .A1(reg_mem[1474]), .A2(n4005), .B1(n6972), .B2(data_w[2]), 
        .ZN(n4007) );
  INV_X1 U2786 ( .A(n4008), .ZN(n6967) );
  AOI22_X1 U2787 ( .A1(reg_mem[1475]), .A2(n4005), .B1(n6972), .B2(data_w[3]), 
        .ZN(n4008) );
  INV_X1 U2788 ( .A(n4009), .ZN(n6968) );
  AOI22_X1 U2789 ( .A1(reg_mem[1476]), .A2(n4005), .B1(n6972), .B2(data_w[4]), 
        .ZN(n4009) );
  INV_X1 U2790 ( .A(n4010), .ZN(n6969) );
  AOI22_X1 U2791 ( .A1(reg_mem[1477]), .A2(n4005), .B1(n6972), .B2(data_w[5]), 
        .ZN(n4010) );
  INV_X1 U2792 ( .A(n4011), .ZN(n6970) );
  AOI22_X1 U2793 ( .A1(reg_mem[1478]), .A2(n4005), .B1(n6972), .B2(data_w[6]), 
        .ZN(n4011) );
  INV_X1 U2794 ( .A(n4012), .ZN(n6971) );
  AOI22_X1 U2795 ( .A1(reg_mem[1479]), .A2(n4005), .B1(n6972), .B2(data_w[7]), 
        .ZN(n4012) );
  INV_X1 U2796 ( .A(n4013), .ZN(n8693) );
  AOI22_X1 U2797 ( .A1(reg_mem[1480]), .A2(n4014), .B1(n8701), .B2(data_w[0]), 
        .ZN(n4013) );
  INV_X1 U2798 ( .A(n4015), .ZN(n8694) );
  AOI22_X1 U2799 ( .A1(reg_mem[1481]), .A2(n4014), .B1(n8701), .B2(data_w[1]), 
        .ZN(n4015) );
  INV_X1 U2800 ( .A(n4016), .ZN(n8695) );
  AOI22_X1 U2801 ( .A1(reg_mem[1482]), .A2(n4014), .B1(n8701), .B2(data_w[2]), 
        .ZN(n4016) );
  INV_X1 U2802 ( .A(n4017), .ZN(n8696) );
  AOI22_X1 U2803 ( .A1(reg_mem[1483]), .A2(n4014), .B1(n8701), .B2(data_w[3]), 
        .ZN(n4017) );
  INV_X1 U2804 ( .A(n4018), .ZN(n8697) );
  AOI22_X1 U2805 ( .A1(reg_mem[1484]), .A2(n4014), .B1(n8701), .B2(data_w[4]), 
        .ZN(n4018) );
  INV_X1 U2806 ( .A(n4019), .ZN(n8698) );
  AOI22_X1 U2807 ( .A1(reg_mem[1485]), .A2(n4014), .B1(n8701), .B2(data_w[5]), 
        .ZN(n4019) );
  INV_X1 U2808 ( .A(n4020), .ZN(n8699) );
  AOI22_X1 U2809 ( .A1(reg_mem[1486]), .A2(n4014), .B1(n8701), .B2(data_w[6]), 
        .ZN(n4020) );
  INV_X1 U2810 ( .A(n4021), .ZN(n8700) );
  AOI22_X1 U2811 ( .A1(reg_mem[1487]), .A2(n4014), .B1(n8701), .B2(data_w[7]), 
        .ZN(n4021) );
  INV_X1 U2812 ( .A(n4022), .ZN(n7540) );
  AOI22_X1 U2813 ( .A1(reg_mem[1488]), .A2(n4023), .B1(n7548), .B2(data_w[0]), 
        .ZN(n4022) );
  INV_X1 U2814 ( .A(n4024), .ZN(n7541) );
  AOI22_X1 U2815 ( .A1(reg_mem[1489]), .A2(n4023), .B1(n7548), .B2(data_w[1]), 
        .ZN(n4024) );
  INV_X1 U2816 ( .A(n4025), .ZN(n7542) );
  AOI22_X1 U2817 ( .A1(reg_mem[1490]), .A2(n4023), .B1(n7548), .B2(data_w[2]), 
        .ZN(n4025) );
  INV_X1 U2818 ( .A(n4026), .ZN(n7543) );
  AOI22_X1 U2819 ( .A1(reg_mem[1491]), .A2(n4023), .B1(n7548), .B2(data_w[3]), 
        .ZN(n4026) );
  INV_X1 U2820 ( .A(n4027), .ZN(n7544) );
  AOI22_X1 U2821 ( .A1(reg_mem[1492]), .A2(n4023), .B1(n7548), .B2(data_w[4]), 
        .ZN(n4027) );
  INV_X1 U2822 ( .A(n4028), .ZN(n7545) );
  AOI22_X1 U2823 ( .A1(reg_mem[1493]), .A2(n4023), .B1(n7548), .B2(data_w[5]), 
        .ZN(n4028) );
  INV_X1 U2824 ( .A(n4029), .ZN(n7546) );
  AOI22_X1 U2825 ( .A1(reg_mem[1494]), .A2(n4023), .B1(n7548), .B2(data_w[6]), 
        .ZN(n4029) );
  INV_X1 U2826 ( .A(n4030), .ZN(n7547) );
  AOI22_X1 U2827 ( .A1(reg_mem[1495]), .A2(n4023), .B1(n7548), .B2(data_w[7]), 
        .ZN(n4030) );
  INV_X1 U2828 ( .A(n4031), .ZN(n8117) );
  AOI22_X1 U2829 ( .A1(reg_mem[1496]), .A2(n4032), .B1(n8125), .B2(data_w[0]), 
        .ZN(n4031) );
  INV_X1 U2830 ( .A(n4033), .ZN(n8118) );
  AOI22_X1 U2831 ( .A1(reg_mem[1497]), .A2(n4032), .B1(n8125), .B2(data_w[1]), 
        .ZN(n4033) );
  INV_X1 U2832 ( .A(n4034), .ZN(n8119) );
  AOI22_X1 U2833 ( .A1(reg_mem[1498]), .A2(n4032), .B1(n8125), .B2(data_w[2]), 
        .ZN(n4034) );
  INV_X1 U2834 ( .A(n4035), .ZN(n8120) );
  AOI22_X1 U2835 ( .A1(reg_mem[1499]), .A2(n4032), .B1(n8125), .B2(data_w[3]), 
        .ZN(n4035) );
  INV_X1 U2836 ( .A(n4036), .ZN(n8121) );
  AOI22_X1 U2837 ( .A1(reg_mem[1500]), .A2(n4032), .B1(n8125), .B2(data_w[4]), 
        .ZN(n4036) );
  INV_X1 U2838 ( .A(n4037), .ZN(n8122) );
  AOI22_X1 U2839 ( .A1(reg_mem[1501]), .A2(n4032), .B1(n8125), .B2(data_w[5]), 
        .ZN(n4037) );
  INV_X1 U2840 ( .A(n4038), .ZN(n8123) );
  AOI22_X1 U2841 ( .A1(reg_mem[1502]), .A2(n4032), .B1(n8125), .B2(data_w[6]), 
        .ZN(n4038) );
  INV_X1 U2842 ( .A(n4039), .ZN(n8124) );
  AOI22_X1 U2843 ( .A1(reg_mem[1503]), .A2(n4032), .B1(n8125), .B2(data_w[7]), 
        .ZN(n4039) );
  INV_X1 U2844 ( .A(n4040), .ZN(n6820) );
  AOI22_X1 U2845 ( .A1(reg_mem[1504]), .A2(n4041), .B1(n6828), .B2(data_w[0]), 
        .ZN(n4040) );
  INV_X1 U2846 ( .A(n4042), .ZN(n6821) );
  AOI22_X1 U2847 ( .A1(reg_mem[1505]), .A2(n4041), .B1(n6828), .B2(data_w[1]), 
        .ZN(n4042) );
  INV_X1 U2848 ( .A(n4043), .ZN(n6822) );
  AOI22_X1 U2849 ( .A1(reg_mem[1506]), .A2(n4041), .B1(n6828), .B2(data_w[2]), 
        .ZN(n4043) );
  INV_X1 U2850 ( .A(n4044), .ZN(n6823) );
  AOI22_X1 U2851 ( .A1(reg_mem[1507]), .A2(n4041), .B1(n6828), .B2(data_w[3]), 
        .ZN(n4044) );
  INV_X1 U2852 ( .A(n4045), .ZN(n6824) );
  AOI22_X1 U2853 ( .A1(reg_mem[1508]), .A2(n4041), .B1(n6828), .B2(data_w[4]), 
        .ZN(n4045) );
  INV_X1 U2854 ( .A(n4046), .ZN(n6825) );
  AOI22_X1 U2855 ( .A1(reg_mem[1509]), .A2(n4041), .B1(n6828), .B2(data_w[5]), 
        .ZN(n4046) );
  INV_X1 U2856 ( .A(n4047), .ZN(n6826) );
  AOI22_X1 U2857 ( .A1(reg_mem[1510]), .A2(n4041), .B1(n6828), .B2(data_w[6]), 
        .ZN(n4047) );
  INV_X1 U2858 ( .A(n4048), .ZN(n6827) );
  AOI22_X1 U2859 ( .A1(reg_mem[1511]), .A2(n4041), .B1(n6828), .B2(data_w[7]), 
        .ZN(n4048) );
  INV_X1 U2860 ( .A(n4049), .ZN(n8549) );
  AOI22_X1 U2861 ( .A1(reg_mem[1512]), .A2(n4050), .B1(n8557), .B2(data_w[0]), 
        .ZN(n4049) );
  INV_X1 U2862 ( .A(n4051), .ZN(n8550) );
  AOI22_X1 U2863 ( .A1(reg_mem[1513]), .A2(n4050), .B1(n8557), .B2(data_w[1]), 
        .ZN(n4051) );
  INV_X1 U2864 ( .A(n4052), .ZN(n8551) );
  AOI22_X1 U2865 ( .A1(reg_mem[1514]), .A2(n4050), .B1(n8557), .B2(data_w[2]), 
        .ZN(n4052) );
  INV_X1 U2866 ( .A(n4053), .ZN(n8552) );
  AOI22_X1 U2867 ( .A1(reg_mem[1515]), .A2(n4050), .B1(n8557), .B2(data_w[3]), 
        .ZN(n4053) );
  INV_X1 U2868 ( .A(n4054), .ZN(n8553) );
  AOI22_X1 U2869 ( .A1(reg_mem[1516]), .A2(n4050), .B1(n8557), .B2(data_w[4]), 
        .ZN(n4054) );
  INV_X1 U2870 ( .A(n4055), .ZN(n8554) );
  AOI22_X1 U2871 ( .A1(reg_mem[1517]), .A2(n4050), .B1(n8557), .B2(data_w[5]), 
        .ZN(n4055) );
  INV_X1 U2872 ( .A(n4056), .ZN(n8555) );
  AOI22_X1 U2873 ( .A1(reg_mem[1518]), .A2(n4050), .B1(n8557), .B2(data_w[6]), 
        .ZN(n4056) );
  INV_X1 U2874 ( .A(n4057), .ZN(n8556) );
  AOI22_X1 U2875 ( .A1(reg_mem[1519]), .A2(n4050), .B1(n8557), .B2(data_w[7]), 
        .ZN(n4057) );
  INV_X1 U2876 ( .A(n4058), .ZN(n7396) );
  AOI22_X1 U2877 ( .A1(reg_mem[1520]), .A2(n4059), .B1(n7404), .B2(data_w[0]), 
        .ZN(n4058) );
  INV_X1 U2878 ( .A(n4060), .ZN(n7397) );
  AOI22_X1 U2879 ( .A1(reg_mem[1521]), .A2(n4059), .B1(n7404), .B2(data_w[1]), 
        .ZN(n4060) );
  INV_X1 U2880 ( .A(n4061), .ZN(n7398) );
  AOI22_X1 U2881 ( .A1(reg_mem[1522]), .A2(n4059), .B1(n7404), .B2(data_w[2]), 
        .ZN(n4061) );
  INV_X1 U2882 ( .A(n4062), .ZN(n7399) );
  AOI22_X1 U2883 ( .A1(reg_mem[1523]), .A2(n4059), .B1(n7404), .B2(data_w[3]), 
        .ZN(n4062) );
  INV_X1 U2884 ( .A(n4063), .ZN(n7400) );
  AOI22_X1 U2885 ( .A1(reg_mem[1524]), .A2(n4059), .B1(n7404), .B2(data_w[4]), 
        .ZN(n4063) );
  INV_X1 U2886 ( .A(n4064), .ZN(n7401) );
  AOI22_X1 U2887 ( .A1(reg_mem[1525]), .A2(n4059), .B1(n7404), .B2(data_w[5]), 
        .ZN(n4064) );
  INV_X1 U2888 ( .A(n4065), .ZN(n7402) );
  AOI22_X1 U2889 ( .A1(reg_mem[1526]), .A2(n4059), .B1(n7404), .B2(data_w[6]), 
        .ZN(n4065) );
  INV_X1 U2890 ( .A(n4066), .ZN(n7403) );
  AOI22_X1 U2891 ( .A1(reg_mem[1527]), .A2(n4059), .B1(n7404), .B2(data_w[7]), 
        .ZN(n4066) );
  INV_X1 U2892 ( .A(n4067), .ZN(n7973) );
  AOI22_X1 U2893 ( .A1(reg_mem[1528]), .A2(n4068), .B1(n7981), .B2(data_w[0]), 
        .ZN(n4067) );
  INV_X1 U2894 ( .A(n4069), .ZN(n7974) );
  AOI22_X1 U2895 ( .A1(reg_mem[1529]), .A2(n4068), .B1(n7981), .B2(data_w[1]), 
        .ZN(n4069) );
  INV_X1 U2896 ( .A(n4070), .ZN(n7975) );
  AOI22_X1 U2897 ( .A1(reg_mem[1530]), .A2(n4068), .B1(n7981), .B2(data_w[2]), 
        .ZN(n4070) );
  INV_X1 U2898 ( .A(n4071), .ZN(n7976) );
  AOI22_X1 U2899 ( .A1(reg_mem[1531]), .A2(n4068), .B1(n7981), .B2(data_w[3]), 
        .ZN(n4071) );
  INV_X1 U2900 ( .A(n4072), .ZN(n7977) );
  AOI22_X1 U2901 ( .A1(reg_mem[1532]), .A2(n4068), .B1(n7981), .B2(data_w[4]), 
        .ZN(n4072) );
  INV_X1 U2902 ( .A(n4073), .ZN(n7978) );
  AOI22_X1 U2903 ( .A1(reg_mem[1533]), .A2(n4068), .B1(n7981), .B2(data_w[5]), 
        .ZN(n4073) );
  INV_X1 U2904 ( .A(n4074), .ZN(n7979) );
  AOI22_X1 U2905 ( .A1(reg_mem[1534]), .A2(n4068), .B1(n7981), .B2(data_w[6]), 
        .ZN(n4074) );
  INV_X1 U2906 ( .A(n4075), .ZN(n7980) );
  AOI22_X1 U2907 ( .A1(reg_mem[1535]), .A2(n4068), .B1(n7981), .B2(data_w[7]), 
        .ZN(n4075) );
  INV_X1 U2908 ( .A(n4076), .ZN(n7243) );
  AOI22_X1 U2909 ( .A1(reg_mem[1536]), .A2(n4077), .B1(n7251), .B2(data_w[0]), 
        .ZN(n4076) );
  INV_X1 U2910 ( .A(n4078), .ZN(n7244) );
  AOI22_X1 U2911 ( .A1(reg_mem[1537]), .A2(n4077), .B1(n7251), .B2(data_w[1]), 
        .ZN(n4078) );
  INV_X1 U2912 ( .A(n4079), .ZN(n7245) );
  AOI22_X1 U2913 ( .A1(reg_mem[1538]), .A2(n4077), .B1(n7251), .B2(data_w[2]), 
        .ZN(n4079) );
  INV_X1 U2914 ( .A(n4080), .ZN(n7246) );
  AOI22_X1 U2915 ( .A1(reg_mem[1539]), .A2(n4077), .B1(n7251), .B2(data_w[3]), 
        .ZN(n4080) );
  INV_X1 U2916 ( .A(n4081), .ZN(n7247) );
  AOI22_X1 U2917 ( .A1(reg_mem[1540]), .A2(n4077), .B1(n7251), .B2(data_w[4]), 
        .ZN(n4081) );
  INV_X1 U2918 ( .A(n4082), .ZN(n7248) );
  AOI22_X1 U2919 ( .A1(reg_mem[1541]), .A2(n4077), .B1(n7251), .B2(data_w[5]), 
        .ZN(n4082) );
  INV_X1 U2920 ( .A(n4083), .ZN(n7249) );
  AOI22_X1 U2921 ( .A1(reg_mem[1542]), .A2(n4077), .B1(n7251), .B2(data_w[6]), 
        .ZN(n4083) );
  INV_X1 U2922 ( .A(n4084), .ZN(n7250) );
  AOI22_X1 U2923 ( .A1(reg_mem[1543]), .A2(n4077), .B1(n7251), .B2(data_w[7]), 
        .ZN(n4084) );
  INV_X1 U2924 ( .A(n4086), .ZN(n8972) );
  AOI22_X1 U2925 ( .A1(reg_mem[1544]), .A2(n4087), .B1(n8980), .B2(data_w[0]), 
        .ZN(n4086) );
  INV_X1 U2926 ( .A(n4088), .ZN(n8973) );
  AOI22_X1 U2927 ( .A1(reg_mem[1545]), .A2(n4087), .B1(n8980), .B2(data_w[1]), 
        .ZN(n4088) );
  INV_X1 U2928 ( .A(n4089), .ZN(n8974) );
  AOI22_X1 U2929 ( .A1(reg_mem[1546]), .A2(n4087), .B1(n8980), .B2(data_w[2]), 
        .ZN(n4089) );
  INV_X1 U2930 ( .A(n4090), .ZN(n8975) );
  AOI22_X1 U2931 ( .A1(reg_mem[1547]), .A2(n4087), .B1(n8980), .B2(data_w[3]), 
        .ZN(n4090) );
  INV_X1 U2932 ( .A(n4091), .ZN(n8976) );
  AOI22_X1 U2933 ( .A1(reg_mem[1548]), .A2(n4087), .B1(n8980), .B2(data_w[4]), 
        .ZN(n4091) );
  INV_X1 U2934 ( .A(n4092), .ZN(n8977) );
  AOI22_X1 U2935 ( .A1(reg_mem[1549]), .A2(n4087), .B1(n8980), .B2(data_w[5]), 
        .ZN(n4092) );
  INV_X1 U2936 ( .A(n4093), .ZN(n8978) );
  AOI22_X1 U2937 ( .A1(reg_mem[1550]), .A2(n4087), .B1(n8980), .B2(data_w[6]), 
        .ZN(n4093) );
  INV_X1 U2938 ( .A(n4094), .ZN(n8979) );
  AOI22_X1 U2939 ( .A1(reg_mem[1551]), .A2(n4087), .B1(n8980), .B2(data_w[7]), 
        .ZN(n4094) );
  INV_X1 U2940 ( .A(n4095), .ZN(n7819) );
  AOI22_X1 U2941 ( .A1(reg_mem[1552]), .A2(n4096), .B1(n7827), .B2(data_w[0]), 
        .ZN(n4095) );
  INV_X1 U2942 ( .A(n4097), .ZN(n7820) );
  AOI22_X1 U2943 ( .A1(reg_mem[1553]), .A2(n4096), .B1(n7827), .B2(data_w[1]), 
        .ZN(n4097) );
  INV_X1 U2944 ( .A(n4098), .ZN(n7821) );
  AOI22_X1 U2945 ( .A1(reg_mem[1554]), .A2(n4096), .B1(n7827), .B2(data_w[2]), 
        .ZN(n4098) );
  INV_X1 U2946 ( .A(n4099), .ZN(n7822) );
  AOI22_X1 U2947 ( .A1(reg_mem[1555]), .A2(n4096), .B1(n7827), .B2(data_w[3]), 
        .ZN(n4099) );
  INV_X1 U2948 ( .A(n4100), .ZN(n7823) );
  AOI22_X1 U2949 ( .A1(reg_mem[1556]), .A2(n4096), .B1(n7827), .B2(data_w[4]), 
        .ZN(n4100) );
  INV_X1 U2950 ( .A(n4101), .ZN(n7824) );
  AOI22_X1 U2951 ( .A1(reg_mem[1557]), .A2(n4096), .B1(n7827), .B2(data_w[5]), 
        .ZN(n4101) );
  INV_X1 U2952 ( .A(n4102), .ZN(n7825) );
  AOI22_X1 U2953 ( .A1(reg_mem[1558]), .A2(n4096), .B1(n7827), .B2(data_w[6]), 
        .ZN(n4102) );
  INV_X1 U2954 ( .A(n4103), .ZN(n7826) );
  AOI22_X1 U2955 ( .A1(reg_mem[1559]), .A2(n4096), .B1(n7827), .B2(data_w[7]), 
        .ZN(n4103) );
  INV_X1 U2956 ( .A(n4104), .ZN(n8396) );
  AOI22_X1 U2957 ( .A1(reg_mem[1560]), .A2(n4105), .B1(n8404), .B2(data_w[0]), 
        .ZN(n4104) );
  INV_X1 U2958 ( .A(n4106), .ZN(n8397) );
  AOI22_X1 U2959 ( .A1(reg_mem[1561]), .A2(n4105), .B1(n8404), .B2(data_w[1]), 
        .ZN(n4106) );
  INV_X1 U2960 ( .A(n4107), .ZN(n8398) );
  AOI22_X1 U2961 ( .A1(reg_mem[1562]), .A2(n4105), .B1(n8404), .B2(data_w[2]), 
        .ZN(n4107) );
  INV_X1 U2962 ( .A(n4108), .ZN(n8399) );
  AOI22_X1 U2963 ( .A1(reg_mem[1563]), .A2(n4105), .B1(n8404), .B2(data_w[3]), 
        .ZN(n4108) );
  INV_X1 U2964 ( .A(n4109), .ZN(n8400) );
  AOI22_X1 U2965 ( .A1(reg_mem[1564]), .A2(n4105), .B1(n8404), .B2(data_w[4]), 
        .ZN(n4109) );
  INV_X1 U2966 ( .A(n4110), .ZN(n8401) );
  AOI22_X1 U2967 ( .A1(reg_mem[1565]), .A2(n4105), .B1(n8404), .B2(data_w[5]), 
        .ZN(n4110) );
  INV_X1 U2968 ( .A(n4111), .ZN(n8402) );
  AOI22_X1 U2969 ( .A1(reg_mem[1566]), .A2(n4105), .B1(n8404), .B2(data_w[6]), 
        .ZN(n4111) );
  INV_X1 U2970 ( .A(n4112), .ZN(n8403) );
  AOI22_X1 U2971 ( .A1(reg_mem[1567]), .A2(n4105), .B1(n8404), .B2(data_w[7]), 
        .ZN(n4112) );
  INV_X1 U2972 ( .A(n4113), .ZN(n7099) );
  AOI22_X1 U2973 ( .A1(reg_mem[1568]), .A2(n4114), .B1(n7107), .B2(data_w[0]), 
        .ZN(n4113) );
  INV_X1 U2974 ( .A(n4115), .ZN(n7100) );
  AOI22_X1 U2975 ( .A1(reg_mem[1569]), .A2(n4114), .B1(n7107), .B2(data_w[1]), 
        .ZN(n4115) );
  INV_X1 U2976 ( .A(n4116), .ZN(n7101) );
  AOI22_X1 U2977 ( .A1(reg_mem[1570]), .A2(n4114), .B1(n7107), .B2(data_w[2]), 
        .ZN(n4116) );
  INV_X1 U2978 ( .A(n4117), .ZN(n7102) );
  AOI22_X1 U2979 ( .A1(reg_mem[1571]), .A2(n4114), .B1(n7107), .B2(data_w[3]), 
        .ZN(n4117) );
  INV_X1 U2980 ( .A(n4118), .ZN(n7103) );
  AOI22_X1 U2981 ( .A1(reg_mem[1572]), .A2(n4114), .B1(n7107), .B2(data_w[4]), 
        .ZN(n4118) );
  INV_X1 U2982 ( .A(n4119), .ZN(n7104) );
  AOI22_X1 U2983 ( .A1(reg_mem[1573]), .A2(n4114), .B1(n7107), .B2(data_w[5]), 
        .ZN(n4119) );
  INV_X1 U2984 ( .A(n4120), .ZN(n7105) );
  AOI22_X1 U2985 ( .A1(reg_mem[1574]), .A2(n4114), .B1(n7107), .B2(data_w[6]), 
        .ZN(n4120) );
  INV_X1 U2986 ( .A(n4121), .ZN(n7106) );
  AOI22_X1 U2987 ( .A1(reg_mem[1575]), .A2(n4114), .B1(n7107), .B2(data_w[7]), 
        .ZN(n4121) );
  INV_X1 U2988 ( .A(n4122), .ZN(n8828) );
  AOI22_X1 U2989 ( .A1(reg_mem[1576]), .A2(n4123), .B1(n8836), .B2(data_w[0]), 
        .ZN(n4122) );
  INV_X1 U2990 ( .A(n4124), .ZN(n8829) );
  AOI22_X1 U2991 ( .A1(reg_mem[1577]), .A2(n4123), .B1(n8836), .B2(data_w[1]), 
        .ZN(n4124) );
  INV_X1 U2992 ( .A(n4125), .ZN(n8830) );
  AOI22_X1 U2993 ( .A1(reg_mem[1578]), .A2(n4123), .B1(n8836), .B2(data_w[2]), 
        .ZN(n4125) );
  INV_X1 U2994 ( .A(n4126), .ZN(n8831) );
  AOI22_X1 U2995 ( .A1(reg_mem[1579]), .A2(n4123), .B1(n8836), .B2(data_w[3]), 
        .ZN(n4126) );
  INV_X1 U2996 ( .A(n4127), .ZN(n8832) );
  AOI22_X1 U2997 ( .A1(reg_mem[1580]), .A2(n4123), .B1(n8836), .B2(data_w[4]), 
        .ZN(n4127) );
  INV_X1 U2998 ( .A(n4128), .ZN(n8833) );
  AOI22_X1 U2999 ( .A1(reg_mem[1581]), .A2(n4123), .B1(n8836), .B2(data_w[5]), 
        .ZN(n4128) );
  INV_X1 U3000 ( .A(n4129), .ZN(n8834) );
  AOI22_X1 U3001 ( .A1(reg_mem[1582]), .A2(n4123), .B1(n8836), .B2(data_w[6]), 
        .ZN(n4129) );
  INV_X1 U3002 ( .A(n4130), .ZN(n8835) );
  AOI22_X1 U3003 ( .A1(reg_mem[1583]), .A2(n4123), .B1(n8836), .B2(data_w[7]), 
        .ZN(n4130) );
  INV_X1 U3004 ( .A(n4131), .ZN(n7675) );
  AOI22_X1 U3005 ( .A1(reg_mem[1584]), .A2(n4132), .B1(n7683), .B2(data_w[0]), 
        .ZN(n4131) );
  INV_X1 U3006 ( .A(n4133), .ZN(n7676) );
  AOI22_X1 U3007 ( .A1(reg_mem[1585]), .A2(n4132), .B1(n7683), .B2(data_w[1]), 
        .ZN(n4133) );
  INV_X1 U3008 ( .A(n4134), .ZN(n7677) );
  AOI22_X1 U3009 ( .A1(reg_mem[1586]), .A2(n4132), .B1(n7683), .B2(data_w[2]), 
        .ZN(n4134) );
  INV_X1 U3010 ( .A(n4135), .ZN(n7678) );
  AOI22_X1 U3011 ( .A1(reg_mem[1587]), .A2(n4132), .B1(n7683), .B2(data_w[3]), 
        .ZN(n4135) );
  INV_X1 U3012 ( .A(n4136), .ZN(n7679) );
  AOI22_X1 U3013 ( .A1(reg_mem[1588]), .A2(n4132), .B1(n7683), .B2(data_w[4]), 
        .ZN(n4136) );
  INV_X1 U3014 ( .A(n4137), .ZN(n7680) );
  AOI22_X1 U3015 ( .A1(reg_mem[1589]), .A2(n4132), .B1(n7683), .B2(data_w[5]), 
        .ZN(n4137) );
  INV_X1 U3016 ( .A(n4138), .ZN(n7681) );
  AOI22_X1 U3017 ( .A1(reg_mem[1590]), .A2(n4132), .B1(n7683), .B2(data_w[6]), 
        .ZN(n4138) );
  INV_X1 U3018 ( .A(n4139), .ZN(n7682) );
  AOI22_X1 U3019 ( .A1(reg_mem[1591]), .A2(n4132), .B1(n7683), .B2(data_w[7]), 
        .ZN(n4139) );
  INV_X1 U3020 ( .A(n4140), .ZN(n8252) );
  AOI22_X1 U3021 ( .A1(reg_mem[1592]), .A2(n4141), .B1(n8260), .B2(data_w[0]), 
        .ZN(n4140) );
  INV_X1 U3022 ( .A(n4142), .ZN(n8253) );
  AOI22_X1 U3023 ( .A1(reg_mem[1593]), .A2(n4141), .B1(n8260), .B2(data_w[1]), 
        .ZN(n4142) );
  INV_X1 U3024 ( .A(n4143), .ZN(n8254) );
  AOI22_X1 U3025 ( .A1(reg_mem[1594]), .A2(n4141), .B1(n8260), .B2(data_w[2]), 
        .ZN(n4143) );
  INV_X1 U3026 ( .A(n4144), .ZN(n8255) );
  AOI22_X1 U3027 ( .A1(reg_mem[1595]), .A2(n4141), .B1(n8260), .B2(data_w[3]), 
        .ZN(n4144) );
  INV_X1 U3028 ( .A(n4145), .ZN(n8256) );
  AOI22_X1 U3029 ( .A1(reg_mem[1596]), .A2(n4141), .B1(n8260), .B2(data_w[4]), 
        .ZN(n4145) );
  INV_X1 U3030 ( .A(n4146), .ZN(n8257) );
  AOI22_X1 U3031 ( .A1(reg_mem[1597]), .A2(n4141), .B1(n8260), .B2(data_w[5]), 
        .ZN(n4146) );
  INV_X1 U3032 ( .A(n4147), .ZN(n8258) );
  AOI22_X1 U3033 ( .A1(reg_mem[1598]), .A2(n4141), .B1(n8260), .B2(data_w[6]), 
        .ZN(n4147) );
  INV_X1 U3034 ( .A(n4148), .ZN(n8259) );
  AOI22_X1 U3035 ( .A1(reg_mem[1599]), .A2(n4141), .B1(n8260), .B2(data_w[7]), 
        .ZN(n4148) );
  INV_X1 U3036 ( .A(n4149), .ZN(n6955) );
  AOI22_X1 U3037 ( .A1(reg_mem[1600]), .A2(n4150), .B1(n6963), .B2(data_w[0]), 
        .ZN(n4149) );
  INV_X1 U3038 ( .A(n4151), .ZN(n6956) );
  AOI22_X1 U3039 ( .A1(reg_mem[1601]), .A2(n4150), .B1(n6963), .B2(data_w[1]), 
        .ZN(n4151) );
  INV_X1 U3040 ( .A(n4152), .ZN(n6957) );
  AOI22_X1 U3041 ( .A1(reg_mem[1602]), .A2(n4150), .B1(n6963), .B2(data_w[2]), 
        .ZN(n4152) );
  INV_X1 U3042 ( .A(n4153), .ZN(n6958) );
  AOI22_X1 U3043 ( .A1(reg_mem[1603]), .A2(n4150), .B1(n6963), .B2(data_w[3]), 
        .ZN(n4153) );
  INV_X1 U3044 ( .A(n4154), .ZN(n6959) );
  AOI22_X1 U3045 ( .A1(reg_mem[1604]), .A2(n4150), .B1(n6963), .B2(data_w[4]), 
        .ZN(n4154) );
  INV_X1 U3046 ( .A(n4155), .ZN(n6960) );
  AOI22_X1 U3047 ( .A1(reg_mem[1605]), .A2(n4150), .B1(n6963), .B2(data_w[5]), 
        .ZN(n4155) );
  INV_X1 U3048 ( .A(n4156), .ZN(n6961) );
  AOI22_X1 U3049 ( .A1(reg_mem[1606]), .A2(n4150), .B1(n6963), .B2(data_w[6]), 
        .ZN(n4156) );
  INV_X1 U3050 ( .A(n4157), .ZN(n6962) );
  AOI22_X1 U3051 ( .A1(reg_mem[1607]), .A2(n4150), .B1(n6963), .B2(data_w[7]), 
        .ZN(n4157) );
  INV_X1 U3052 ( .A(n4158), .ZN(n8684) );
  AOI22_X1 U3053 ( .A1(reg_mem[1608]), .A2(n4159), .B1(n8692), .B2(data_w[0]), 
        .ZN(n4158) );
  INV_X1 U3054 ( .A(n4160), .ZN(n8685) );
  AOI22_X1 U3055 ( .A1(reg_mem[1609]), .A2(n4159), .B1(n8692), .B2(data_w[1]), 
        .ZN(n4160) );
  INV_X1 U3056 ( .A(n4161), .ZN(n8686) );
  AOI22_X1 U3057 ( .A1(reg_mem[1610]), .A2(n4159), .B1(n8692), .B2(data_w[2]), 
        .ZN(n4161) );
  INV_X1 U3058 ( .A(n4162), .ZN(n8687) );
  AOI22_X1 U3059 ( .A1(reg_mem[1611]), .A2(n4159), .B1(n8692), .B2(data_w[3]), 
        .ZN(n4162) );
  INV_X1 U3060 ( .A(n4163), .ZN(n8688) );
  AOI22_X1 U3061 ( .A1(reg_mem[1612]), .A2(n4159), .B1(n8692), .B2(data_w[4]), 
        .ZN(n4163) );
  INV_X1 U3062 ( .A(n4164), .ZN(n8689) );
  AOI22_X1 U3063 ( .A1(reg_mem[1613]), .A2(n4159), .B1(n8692), .B2(data_w[5]), 
        .ZN(n4164) );
  INV_X1 U3064 ( .A(n4165), .ZN(n8690) );
  AOI22_X1 U3065 ( .A1(reg_mem[1614]), .A2(n4159), .B1(n8692), .B2(data_w[6]), 
        .ZN(n4165) );
  INV_X1 U3066 ( .A(n4166), .ZN(n8691) );
  AOI22_X1 U3067 ( .A1(reg_mem[1615]), .A2(n4159), .B1(n8692), .B2(data_w[7]), 
        .ZN(n4166) );
  INV_X1 U3068 ( .A(n4167), .ZN(n7531) );
  AOI22_X1 U3069 ( .A1(reg_mem[1616]), .A2(n4168), .B1(n7539), .B2(data_w[0]), 
        .ZN(n4167) );
  INV_X1 U3070 ( .A(n4169), .ZN(n7532) );
  AOI22_X1 U3071 ( .A1(reg_mem[1617]), .A2(n4168), .B1(n7539), .B2(data_w[1]), 
        .ZN(n4169) );
  INV_X1 U3072 ( .A(n4170), .ZN(n7533) );
  AOI22_X1 U3073 ( .A1(reg_mem[1618]), .A2(n4168), .B1(n7539), .B2(data_w[2]), 
        .ZN(n4170) );
  INV_X1 U3074 ( .A(n4171), .ZN(n7534) );
  AOI22_X1 U3075 ( .A1(reg_mem[1619]), .A2(n4168), .B1(n7539), .B2(data_w[3]), 
        .ZN(n4171) );
  INV_X1 U3076 ( .A(n4172), .ZN(n7535) );
  AOI22_X1 U3077 ( .A1(reg_mem[1620]), .A2(n4168), .B1(n7539), .B2(data_w[4]), 
        .ZN(n4172) );
  INV_X1 U3078 ( .A(n4173), .ZN(n7536) );
  AOI22_X1 U3079 ( .A1(reg_mem[1621]), .A2(n4168), .B1(n7539), .B2(data_w[5]), 
        .ZN(n4173) );
  INV_X1 U3080 ( .A(n4174), .ZN(n7537) );
  AOI22_X1 U3081 ( .A1(reg_mem[1622]), .A2(n4168), .B1(n7539), .B2(data_w[6]), 
        .ZN(n4174) );
  INV_X1 U3082 ( .A(n4175), .ZN(n7538) );
  AOI22_X1 U3083 ( .A1(reg_mem[1623]), .A2(n4168), .B1(n7539), .B2(data_w[7]), 
        .ZN(n4175) );
  INV_X1 U3084 ( .A(n4176), .ZN(n8108) );
  AOI22_X1 U3085 ( .A1(reg_mem[1624]), .A2(n4177), .B1(n8116), .B2(data_w[0]), 
        .ZN(n4176) );
  INV_X1 U3086 ( .A(n4178), .ZN(n8109) );
  AOI22_X1 U3087 ( .A1(reg_mem[1625]), .A2(n4177), .B1(n8116), .B2(data_w[1]), 
        .ZN(n4178) );
  INV_X1 U3088 ( .A(n4179), .ZN(n8110) );
  AOI22_X1 U3089 ( .A1(reg_mem[1626]), .A2(n4177), .B1(n8116), .B2(data_w[2]), 
        .ZN(n4179) );
  INV_X1 U3090 ( .A(n4180), .ZN(n8111) );
  AOI22_X1 U3091 ( .A1(reg_mem[1627]), .A2(n4177), .B1(n8116), .B2(data_w[3]), 
        .ZN(n4180) );
  INV_X1 U3092 ( .A(n4181), .ZN(n8112) );
  AOI22_X1 U3093 ( .A1(reg_mem[1628]), .A2(n4177), .B1(n8116), .B2(data_w[4]), 
        .ZN(n4181) );
  INV_X1 U3094 ( .A(n4182), .ZN(n8113) );
  AOI22_X1 U3095 ( .A1(reg_mem[1629]), .A2(n4177), .B1(n8116), .B2(data_w[5]), 
        .ZN(n4182) );
  INV_X1 U3096 ( .A(n4183), .ZN(n8114) );
  AOI22_X1 U3097 ( .A1(reg_mem[1630]), .A2(n4177), .B1(n8116), .B2(data_w[6]), 
        .ZN(n4183) );
  INV_X1 U3098 ( .A(n4184), .ZN(n8115) );
  AOI22_X1 U3099 ( .A1(reg_mem[1631]), .A2(n4177), .B1(n8116), .B2(data_w[7]), 
        .ZN(n4184) );
  INV_X1 U3100 ( .A(n4185), .ZN(n6811) );
  AOI22_X1 U3101 ( .A1(reg_mem[1632]), .A2(n4186), .B1(n6819), .B2(data_w[0]), 
        .ZN(n4185) );
  INV_X1 U3102 ( .A(n4187), .ZN(n6812) );
  AOI22_X1 U3103 ( .A1(reg_mem[1633]), .A2(n4186), .B1(n6819), .B2(data_w[1]), 
        .ZN(n4187) );
  INV_X1 U3104 ( .A(n4188), .ZN(n6813) );
  AOI22_X1 U3105 ( .A1(reg_mem[1634]), .A2(n4186), .B1(n6819), .B2(data_w[2]), 
        .ZN(n4188) );
  INV_X1 U3106 ( .A(n4189), .ZN(n6814) );
  AOI22_X1 U3107 ( .A1(reg_mem[1635]), .A2(n4186), .B1(n6819), .B2(data_w[3]), 
        .ZN(n4189) );
  INV_X1 U3108 ( .A(n4190), .ZN(n6815) );
  AOI22_X1 U3109 ( .A1(reg_mem[1636]), .A2(n4186), .B1(n6819), .B2(data_w[4]), 
        .ZN(n4190) );
  INV_X1 U3110 ( .A(n4191), .ZN(n6816) );
  AOI22_X1 U3111 ( .A1(reg_mem[1637]), .A2(n4186), .B1(n6819), .B2(data_w[5]), 
        .ZN(n4191) );
  INV_X1 U3112 ( .A(n4192), .ZN(n6817) );
  AOI22_X1 U3113 ( .A1(reg_mem[1638]), .A2(n4186), .B1(n6819), .B2(data_w[6]), 
        .ZN(n4192) );
  INV_X1 U3114 ( .A(n4193), .ZN(n6818) );
  AOI22_X1 U3115 ( .A1(reg_mem[1639]), .A2(n4186), .B1(n6819), .B2(data_w[7]), 
        .ZN(n4193) );
  INV_X1 U3116 ( .A(n4194), .ZN(n8540) );
  AOI22_X1 U3117 ( .A1(reg_mem[1640]), .A2(n4195), .B1(n8548), .B2(data_w[0]), 
        .ZN(n4194) );
  INV_X1 U3118 ( .A(n4196), .ZN(n8541) );
  AOI22_X1 U3119 ( .A1(reg_mem[1641]), .A2(n4195), .B1(n8548), .B2(data_w[1]), 
        .ZN(n4196) );
  INV_X1 U3120 ( .A(n4197), .ZN(n8542) );
  AOI22_X1 U3121 ( .A1(reg_mem[1642]), .A2(n4195), .B1(n8548), .B2(data_w[2]), 
        .ZN(n4197) );
  INV_X1 U3122 ( .A(n4198), .ZN(n8543) );
  AOI22_X1 U3123 ( .A1(reg_mem[1643]), .A2(n4195), .B1(n8548), .B2(data_w[3]), 
        .ZN(n4198) );
  INV_X1 U3124 ( .A(n4199), .ZN(n8544) );
  AOI22_X1 U3125 ( .A1(reg_mem[1644]), .A2(n4195), .B1(n8548), .B2(data_w[4]), 
        .ZN(n4199) );
  INV_X1 U3126 ( .A(n4200), .ZN(n8545) );
  AOI22_X1 U3127 ( .A1(reg_mem[1645]), .A2(n4195), .B1(n8548), .B2(data_w[5]), 
        .ZN(n4200) );
  INV_X1 U3128 ( .A(n4201), .ZN(n8546) );
  AOI22_X1 U3129 ( .A1(reg_mem[1646]), .A2(n4195), .B1(n8548), .B2(data_w[6]), 
        .ZN(n4201) );
  INV_X1 U3130 ( .A(n4202), .ZN(n8547) );
  AOI22_X1 U3131 ( .A1(reg_mem[1647]), .A2(n4195), .B1(n8548), .B2(data_w[7]), 
        .ZN(n4202) );
  INV_X1 U3132 ( .A(n4203), .ZN(n7387) );
  AOI22_X1 U3133 ( .A1(reg_mem[1648]), .A2(n4204), .B1(n7395), .B2(data_w[0]), 
        .ZN(n4203) );
  INV_X1 U3134 ( .A(n4205), .ZN(n7388) );
  AOI22_X1 U3135 ( .A1(reg_mem[1649]), .A2(n4204), .B1(n7395), .B2(data_w[1]), 
        .ZN(n4205) );
  INV_X1 U3136 ( .A(n4206), .ZN(n7389) );
  AOI22_X1 U3137 ( .A1(reg_mem[1650]), .A2(n4204), .B1(n7395), .B2(data_w[2]), 
        .ZN(n4206) );
  INV_X1 U3138 ( .A(n4207), .ZN(n7390) );
  AOI22_X1 U3139 ( .A1(reg_mem[1651]), .A2(n4204), .B1(n7395), .B2(data_w[3]), 
        .ZN(n4207) );
  INV_X1 U3140 ( .A(n4208), .ZN(n7391) );
  AOI22_X1 U3141 ( .A1(reg_mem[1652]), .A2(n4204), .B1(n7395), .B2(data_w[4]), 
        .ZN(n4208) );
  INV_X1 U3142 ( .A(n4209), .ZN(n7392) );
  AOI22_X1 U3143 ( .A1(reg_mem[1653]), .A2(n4204), .B1(n7395), .B2(data_w[5]), 
        .ZN(n4209) );
  INV_X1 U3144 ( .A(n4210), .ZN(n7393) );
  AOI22_X1 U3145 ( .A1(reg_mem[1654]), .A2(n4204), .B1(n7395), .B2(data_w[6]), 
        .ZN(n4210) );
  INV_X1 U3146 ( .A(n4211), .ZN(n7394) );
  AOI22_X1 U3147 ( .A1(reg_mem[1655]), .A2(n4204), .B1(n7395), .B2(data_w[7]), 
        .ZN(n4211) );
  INV_X1 U3148 ( .A(n4212), .ZN(n7964) );
  AOI22_X1 U3149 ( .A1(reg_mem[1656]), .A2(n4213), .B1(n7972), .B2(data_w[0]), 
        .ZN(n4212) );
  INV_X1 U3150 ( .A(n4214), .ZN(n7965) );
  AOI22_X1 U3151 ( .A1(reg_mem[1657]), .A2(n4213), .B1(n7972), .B2(data_w[1]), 
        .ZN(n4214) );
  INV_X1 U3152 ( .A(n4215), .ZN(n7966) );
  AOI22_X1 U3153 ( .A1(reg_mem[1658]), .A2(n4213), .B1(n7972), .B2(data_w[2]), 
        .ZN(n4215) );
  INV_X1 U3154 ( .A(n4216), .ZN(n7967) );
  AOI22_X1 U3155 ( .A1(reg_mem[1659]), .A2(n4213), .B1(n7972), .B2(data_w[3]), 
        .ZN(n4216) );
  INV_X1 U3156 ( .A(n4217), .ZN(n7968) );
  AOI22_X1 U3157 ( .A1(reg_mem[1660]), .A2(n4213), .B1(n7972), .B2(data_w[4]), 
        .ZN(n4217) );
  INV_X1 U3158 ( .A(n4218), .ZN(n7969) );
  AOI22_X1 U3159 ( .A1(reg_mem[1661]), .A2(n4213), .B1(n7972), .B2(data_w[5]), 
        .ZN(n4218) );
  INV_X1 U3160 ( .A(n4219), .ZN(n7970) );
  AOI22_X1 U3161 ( .A1(reg_mem[1662]), .A2(n4213), .B1(n7972), .B2(data_w[6]), 
        .ZN(n4219) );
  INV_X1 U3162 ( .A(n4220), .ZN(n7971) );
  AOI22_X1 U3163 ( .A1(reg_mem[1663]), .A2(n4213), .B1(n7972), .B2(data_w[7]), 
        .ZN(n4220) );
  INV_X1 U3164 ( .A(n4222), .ZN(n7234) );
  AOI22_X1 U3165 ( .A1(reg_mem[1664]), .A2(n4223), .B1(n7242), .B2(data_w[0]), 
        .ZN(n4222) );
  INV_X1 U3166 ( .A(n4224), .ZN(n7235) );
  AOI22_X1 U3167 ( .A1(reg_mem[1665]), .A2(n4223), .B1(n7242), .B2(data_w[1]), 
        .ZN(n4224) );
  INV_X1 U3168 ( .A(n4225), .ZN(n7236) );
  AOI22_X1 U3169 ( .A1(reg_mem[1666]), .A2(n4223), .B1(n7242), .B2(data_w[2]), 
        .ZN(n4225) );
  INV_X1 U3170 ( .A(n4226), .ZN(n7237) );
  AOI22_X1 U3171 ( .A1(reg_mem[1667]), .A2(n4223), .B1(n7242), .B2(data_w[3]), 
        .ZN(n4226) );
  INV_X1 U3172 ( .A(n4227), .ZN(n7238) );
  AOI22_X1 U3173 ( .A1(reg_mem[1668]), .A2(n4223), .B1(n7242), .B2(data_w[4]), 
        .ZN(n4227) );
  INV_X1 U3174 ( .A(n4228), .ZN(n7239) );
  AOI22_X1 U3175 ( .A1(reg_mem[1669]), .A2(n4223), .B1(n7242), .B2(data_w[5]), 
        .ZN(n4228) );
  INV_X1 U3176 ( .A(n4229), .ZN(n7240) );
  AOI22_X1 U3177 ( .A1(reg_mem[1670]), .A2(n4223), .B1(n7242), .B2(data_w[6]), 
        .ZN(n4229) );
  INV_X1 U3178 ( .A(n4230), .ZN(n7241) );
  AOI22_X1 U3179 ( .A1(reg_mem[1671]), .A2(n4223), .B1(n7242), .B2(data_w[7]), 
        .ZN(n4230) );
  INV_X1 U3180 ( .A(n4232), .ZN(n8963) );
  AOI22_X1 U3181 ( .A1(reg_mem[1672]), .A2(n4233), .B1(n8971), .B2(data_w[0]), 
        .ZN(n4232) );
  INV_X1 U3182 ( .A(n4234), .ZN(n8964) );
  AOI22_X1 U3183 ( .A1(reg_mem[1673]), .A2(n4233), .B1(n8971), .B2(data_w[1]), 
        .ZN(n4234) );
  INV_X1 U3184 ( .A(n4235), .ZN(n8965) );
  AOI22_X1 U3185 ( .A1(reg_mem[1674]), .A2(n4233), .B1(n8971), .B2(data_w[2]), 
        .ZN(n4235) );
  INV_X1 U3186 ( .A(n4236), .ZN(n8966) );
  AOI22_X1 U3187 ( .A1(reg_mem[1675]), .A2(n4233), .B1(n8971), .B2(data_w[3]), 
        .ZN(n4236) );
  INV_X1 U3188 ( .A(n4237), .ZN(n8967) );
  AOI22_X1 U3189 ( .A1(reg_mem[1676]), .A2(n4233), .B1(n8971), .B2(data_w[4]), 
        .ZN(n4237) );
  INV_X1 U3190 ( .A(n4238), .ZN(n8968) );
  AOI22_X1 U3191 ( .A1(reg_mem[1677]), .A2(n4233), .B1(n8971), .B2(data_w[5]), 
        .ZN(n4238) );
  INV_X1 U3192 ( .A(n4239), .ZN(n8969) );
  AOI22_X1 U3193 ( .A1(reg_mem[1678]), .A2(n4233), .B1(n8971), .B2(data_w[6]), 
        .ZN(n4239) );
  INV_X1 U3194 ( .A(n4240), .ZN(n8970) );
  AOI22_X1 U3195 ( .A1(reg_mem[1679]), .A2(n4233), .B1(n8971), .B2(data_w[7]), 
        .ZN(n4240) );
  INV_X1 U3196 ( .A(n4241), .ZN(n7810) );
  AOI22_X1 U3197 ( .A1(reg_mem[1680]), .A2(n4242), .B1(n7818), .B2(data_w[0]), 
        .ZN(n4241) );
  INV_X1 U3198 ( .A(n4243), .ZN(n7811) );
  AOI22_X1 U3199 ( .A1(reg_mem[1681]), .A2(n4242), .B1(n7818), .B2(data_w[1]), 
        .ZN(n4243) );
  INV_X1 U3200 ( .A(n4244), .ZN(n7812) );
  AOI22_X1 U3201 ( .A1(reg_mem[1682]), .A2(n4242), .B1(n7818), .B2(data_w[2]), 
        .ZN(n4244) );
  INV_X1 U3202 ( .A(n4245), .ZN(n7813) );
  AOI22_X1 U3203 ( .A1(reg_mem[1683]), .A2(n4242), .B1(n7818), .B2(data_w[3]), 
        .ZN(n4245) );
  INV_X1 U3204 ( .A(n4246), .ZN(n7814) );
  AOI22_X1 U3205 ( .A1(reg_mem[1684]), .A2(n4242), .B1(n7818), .B2(data_w[4]), 
        .ZN(n4246) );
  INV_X1 U3206 ( .A(n4247), .ZN(n7815) );
  AOI22_X1 U3207 ( .A1(reg_mem[1685]), .A2(n4242), .B1(n7818), .B2(data_w[5]), 
        .ZN(n4247) );
  INV_X1 U3208 ( .A(n4248), .ZN(n7816) );
  AOI22_X1 U3209 ( .A1(reg_mem[1686]), .A2(n4242), .B1(n7818), .B2(data_w[6]), 
        .ZN(n4248) );
  INV_X1 U3210 ( .A(n4249), .ZN(n7817) );
  AOI22_X1 U3211 ( .A1(reg_mem[1687]), .A2(n4242), .B1(n7818), .B2(data_w[7]), 
        .ZN(n4249) );
  INV_X1 U3212 ( .A(n4250), .ZN(n8387) );
  AOI22_X1 U3213 ( .A1(reg_mem[1688]), .A2(n4251), .B1(n8395), .B2(data_w[0]), 
        .ZN(n4250) );
  INV_X1 U3214 ( .A(n4252), .ZN(n8388) );
  AOI22_X1 U3215 ( .A1(reg_mem[1689]), .A2(n4251), .B1(n8395), .B2(data_w[1]), 
        .ZN(n4252) );
  INV_X1 U3216 ( .A(n4253), .ZN(n8389) );
  AOI22_X1 U3217 ( .A1(reg_mem[1690]), .A2(n4251), .B1(n8395), .B2(data_w[2]), 
        .ZN(n4253) );
  INV_X1 U3218 ( .A(n4254), .ZN(n8390) );
  AOI22_X1 U3219 ( .A1(reg_mem[1691]), .A2(n4251), .B1(n8395), .B2(data_w[3]), 
        .ZN(n4254) );
  INV_X1 U3220 ( .A(n4255), .ZN(n8391) );
  AOI22_X1 U3221 ( .A1(reg_mem[1692]), .A2(n4251), .B1(n8395), .B2(data_w[4]), 
        .ZN(n4255) );
  INV_X1 U3222 ( .A(n4256), .ZN(n8392) );
  AOI22_X1 U3223 ( .A1(reg_mem[1693]), .A2(n4251), .B1(n8395), .B2(data_w[5]), 
        .ZN(n4256) );
  INV_X1 U3224 ( .A(n4257), .ZN(n8393) );
  AOI22_X1 U3225 ( .A1(reg_mem[1694]), .A2(n4251), .B1(n8395), .B2(data_w[6]), 
        .ZN(n4257) );
  INV_X1 U3226 ( .A(n4258), .ZN(n8394) );
  AOI22_X1 U3227 ( .A1(reg_mem[1695]), .A2(n4251), .B1(n8395), .B2(data_w[7]), 
        .ZN(n4258) );
  INV_X1 U3228 ( .A(n4259), .ZN(n7090) );
  AOI22_X1 U3229 ( .A1(reg_mem[1696]), .A2(n4260), .B1(n7098), .B2(data_w[0]), 
        .ZN(n4259) );
  INV_X1 U3230 ( .A(n4261), .ZN(n7091) );
  AOI22_X1 U3231 ( .A1(reg_mem[1697]), .A2(n4260), .B1(n7098), .B2(data_w[1]), 
        .ZN(n4261) );
  INV_X1 U3232 ( .A(n4262), .ZN(n7092) );
  AOI22_X1 U3233 ( .A1(reg_mem[1698]), .A2(n4260), .B1(n7098), .B2(data_w[2]), 
        .ZN(n4262) );
  INV_X1 U3234 ( .A(n4263), .ZN(n7093) );
  AOI22_X1 U3235 ( .A1(reg_mem[1699]), .A2(n4260), .B1(n7098), .B2(data_w[3]), 
        .ZN(n4263) );
  INV_X1 U3236 ( .A(n4264), .ZN(n7094) );
  AOI22_X1 U3237 ( .A1(reg_mem[1700]), .A2(n4260), .B1(n7098), .B2(data_w[4]), 
        .ZN(n4264) );
  INV_X1 U3238 ( .A(n4265), .ZN(n7095) );
  AOI22_X1 U3239 ( .A1(reg_mem[1701]), .A2(n4260), .B1(n7098), .B2(data_w[5]), 
        .ZN(n4265) );
  INV_X1 U3240 ( .A(n4266), .ZN(n7096) );
  AOI22_X1 U3241 ( .A1(reg_mem[1702]), .A2(n4260), .B1(n7098), .B2(data_w[6]), 
        .ZN(n4266) );
  INV_X1 U3242 ( .A(n4267), .ZN(n7097) );
  AOI22_X1 U3243 ( .A1(reg_mem[1703]), .A2(n4260), .B1(n7098), .B2(data_w[7]), 
        .ZN(n4267) );
  INV_X1 U3244 ( .A(n4268), .ZN(n8819) );
  AOI22_X1 U3245 ( .A1(reg_mem[1704]), .A2(n4269), .B1(n8827), .B2(data_w[0]), 
        .ZN(n4268) );
  INV_X1 U3246 ( .A(n4270), .ZN(n8820) );
  AOI22_X1 U3247 ( .A1(reg_mem[1705]), .A2(n4269), .B1(n8827), .B2(data_w[1]), 
        .ZN(n4270) );
  INV_X1 U3248 ( .A(n4271), .ZN(n8821) );
  AOI22_X1 U3249 ( .A1(reg_mem[1706]), .A2(n4269), .B1(n8827), .B2(data_w[2]), 
        .ZN(n4271) );
  INV_X1 U3250 ( .A(n4272), .ZN(n8822) );
  AOI22_X1 U3251 ( .A1(reg_mem[1707]), .A2(n4269), .B1(n8827), .B2(data_w[3]), 
        .ZN(n4272) );
  INV_X1 U3252 ( .A(n4273), .ZN(n8823) );
  AOI22_X1 U3253 ( .A1(reg_mem[1708]), .A2(n4269), .B1(n8827), .B2(data_w[4]), 
        .ZN(n4273) );
  INV_X1 U3254 ( .A(n4274), .ZN(n8824) );
  AOI22_X1 U3255 ( .A1(reg_mem[1709]), .A2(n4269), .B1(n8827), .B2(data_w[5]), 
        .ZN(n4274) );
  INV_X1 U3256 ( .A(n4275), .ZN(n8825) );
  AOI22_X1 U3257 ( .A1(reg_mem[1710]), .A2(n4269), .B1(n8827), .B2(data_w[6]), 
        .ZN(n4275) );
  INV_X1 U3258 ( .A(n4276), .ZN(n8826) );
  AOI22_X1 U3259 ( .A1(reg_mem[1711]), .A2(n4269), .B1(n8827), .B2(data_w[7]), 
        .ZN(n4276) );
  INV_X1 U3260 ( .A(n4277), .ZN(n7666) );
  AOI22_X1 U3261 ( .A1(reg_mem[1712]), .A2(n4278), .B1(n7674), .B2(data_w[0]), 
        .ZN(n4277) );
  INV_X1 U3262 ( .A(n4279), .ZN(n7667) );
  AOI22_X1 U3263 ( .A1(reg_mem[1713]), .A2(n4278), .B1(n7674), .B2(data_w[1]), 
        .ZN(n4279) );
  INV_X1 U3264 ( .A(n4280), .ZN(n7668) );
  AOI22_X1 U3265 ( .A1(reg_mem[1714]), .A2(n4278), .B1(n7674), .B2(data_w[2]), 
        .ZN(n4280) );
  INV_X1 U3266 ( .A(n4281), .ZN(n7669) );
  AOI22_X1 U3267 ( .A1(reg_mem[1715]), .A2(n4278), .B1(n7674), .B2(data_w[3]), 
        .ZN(n4281) );
  INV_X1 U3268 ( .A(n4282), .ZN(n7670) );
  AOI22_X1 U3269 ( .A1(reg_mem[1716]), .A2(n4278), .B1(n7674), .B2(data_w[4]), 
        .ZN(n4282) );
  INV_X1 U3270 ( .A(n4283), .ZN(n7671) );
  AOI22_X1 U3271 ( .A1(reg_mem[1717]), .A2(n4278), .B1(n7674), .B2(data_w[5]), 
        .ZN(n4283) );
  INV_X1 U3272 ( .A(n4284), .ZN(n7672) );
  AOI22_X1 U3273 ( .A1(reg_mem[1718]), .A2(n4278), .B1(n7674), .B2(data_w[6]), 
        .ZN(n4284) );
  INV_X1 U3274 ( .A(n4285), .ZN(n7673) );
  AOI22_X1 U3275 ( .A1(reg_mem[1719]), .A2(n4278), .B1(n7674), .B2(data_w[7]), 
        .ZN(n4285) );
  INV_X1 U3276 ( .A(n4286), .ZN(n8243) );
  AOI22_X1 U3277 ( .A1(reg_mem[1720]), .A2(n4287), .B1(n8251), .B2(data_w[0]), 
        .ZN(n4286) );
  INV_X1 U3278 ( .A(n4288), .ZN(n8244) );
  AOI22_X1 U3279 ( .A1(reg_mem[1721]), .A2(n4287), .B1(n8251), .B2(data_w[1]), 
        .ZN(n4288) );
  INV_X1 U3280 ( .A(n4289), .ZN(n8245) );
  AOI22_X1 U3281 ( .A1(reg_mem[1722]), .A2(n4287), .B1(n8251), .B2(data_w[2]), 
        .ZN(n4289) );
  INV_X1 U3282 ( .A(n4290), .ZN(n8246) );
  AOI22_X1 U3283 ( .A1(reg_mem[1723]), .A2(n4287), .B1(n8251), .B2(data_w[3]), 
        .ZN(n4290) );
  INV_X1 U3284 ( .A(n4291), .ZN(n8247) );
  AOI22_X1 U3285 ( .A1(reg_mem[1724]), .A2(n4287), .B1(n8251), .B2(data_w[4]), 
        .ZN(n4291) );
  INV_X1 U3286 ( .A(n4292), .ZN(n8248) );
  AOI22_X1 U3287 ( .A1(reg_mem[1725]), .A2(n4287), .B1(n8251), .B2(data_w[5]), 
        .ZN(n4292) );
  INV_X1 U3288 ( .A(n4293), .ZN(n8249) );
  AOI22_X1 U3289 ( .A1(reg_mem[1726]), .A2(n4287), .B1(n8251), .B2(data_w[6]), 
        .ZN(n4293) );
  INV_X1 U3290 ( .A(n4294), .ZN(n8250) );
  AOI22_X1 U3291 ( .A1(reg_mem[1727]), .A2(n4287), .B1(n8251), .B2(data_w[7]), 
        .ZN(n4294) );
  INV_X1 U3292 ( .A(n4295), .ZN(n6946) );
  AOI22_X1 U3293 ( .A1(reg_mem[1728]), .A2(n4296), .B1(n6954), .B2(data_w[0]), 
        .ZN(n4295) );
  INV_X1 U3294 ( .A(n4297), .ZN(n6947) );
  AOI22_X1 U3295 ( .A1(reg_mem[1729]), .A2(n4296), .B1(n6954), .B2(data_w[1]), 
        .ZN(n4297) );
  INV_X1 U3296 ( .A(n4298), .ZN(n6948) );
  AOI22_X1 U3297 ( .A1(reg_mem[1730]), .A2(n4296), .B1(n6954), .B2(data_w[2]), 
        .ZN(n4298) );
  INV_X1 U3298 ( .A(n4299), .ZN(n6949) );
  AOI22_X1 U3299 ( .A1(reg_mem[1731]), .A2(n4296), .B1(n6954), .B2(data_w[3]), 
        .ZN(n4299) );
  INV_X1 U3300 ( .A(n4300), .ZN(n6950) );
  AOI22_X1 U3301 ( .A1(reg_mem[1732]), .A2(n4296), .B1(n6954), .B2(data_w[4]), 
        .ZN(n4300) );
  INV_X1 U3302 ( .A(n4301), .ZN(n6951) );
  AOI22_X1 U3303 ( .A1(reg_mem[1733]), .A2(n4296), .B1(n6954), .B2(data_w[5]), 
        .ZN(n4301) );
  INV_X1 U3304 ( .A(n4302), .ZN(n6952) );
  AOI22_X1 U3305 ( .A1(reg_mem[1734]), .A2(n4296), .B1(n6954), .B2(data_w[6]), 
        .ZN(n4302) );
  INV_X1 U3306 ( .A(n4303), .ZN(n6953) );
  AOI22_X1 U3307 ( .A1(reg_mem[1735]), .A2(n4296), .B1(n6954), .B2(data_w[7]), 
        .ZN(n4303) );
  INV_X1 U3308 ( .A(n4304), .ZN(n8675) );
  AOI22_X1 U3309 ( .A1(reg_mem[1736]), .A2(n4305), .B1(n8683), .B2(data_w[0]), 
        .ZN(n4304) );
  INV_X1 U3310 ( .A(n4306), .ZN(n8676) );
  AOI22_X1 U3311 ( .A1(reg_mem[1737]), .A2(n4305), .B1(n8683), .B2(data_w[1]), 
        .ZN(n4306) );
  INV_X1 U3312 ( .A(n4307), .ZN(n8677) );
  AOI22_X1 U3313 ( .A1(reg_mem[1738]), .A2(n4305), .B1(n8683), .B2(data_w[2]), 
        .ZN(n4307) );
  INV_X1 U3314 ( .A(n4308), .ZN(n8678) );
  AOI22_X1 U3315 ( .A1(reg_mem[1739]), .A2(n4305), .B1(n8683), .B2(data_w[3]), 
        .ZN(n4308) );
  INV_X1 U3316 ( .A(n4309), .ZN(n8679) );
  AOI22_X1 U3317 ( .A1(reg_mem[1740]), .A2(n4305), .B1(n8683), .B2(data_w[4]), 
        .ZN(n4309) );
  INV_X1 U3318 ( .A(n4310), .ZN(n8680) );
  AOI22_X1 U3319 ( .A1(reg_mem[1741]), .A2(n4305), .B1(n8683), .B2(data_w[5]), 
        .ZN(n4310) );
  INV_X1 U3320 ( .A(n4311), .ZN(n8681) );
  AOI22_X1 U3321 ( .A1(reg_mem[1742]), .A2(n4305), .B1(n8683), .B2(data_w[6]), 
        .ZN(n4311) );
  INV_X1 U3322 ( .A(n4312), .ZN(n8682) );
  AOI22_X1 U3323 ( .A1(reg_mem[1743]), .A2(n4305), .B1(n8683), .B2(data_w[7]), 
        .ZN(n4312) );
  INV_X1 U3324 ( .A(n4313), .ZN(n7522) );
  AOI22_X1 U3325 ( .A1(reg_mem[1744]), .A2(n4314), .B1(n7530), .B2(data_w[0]), 
        .ZN(n4313) );
  INV_X1 U3326 ( .A(n4315), .ZN(n7523) );
  AOI22_X1 U3327 ( .A1(reg_mem[1745]), .A2(n4314), .B1(n7530), .B2(data_w[1]), 
        .ZN(n4315) );
  INV_X1 U3328 ( .A(n4316), .ZN(n7524) );
  AOI22_X1 U3329 ( .A1(reg_mem[1746]), .A2(n4314), .B1(n7530), .B2(data_w[2]), 
        .ZN(n4316) );
  INV_X1 U3330 ( .A(n4317), .ZN(n7525) );
  AOI22_X1 U3331 ( .A1(reg_mem[1747]), .A2(n4314), .B1(n7530), .B2(data_w[3]), 
        .ZN(n4317) );
  INV_X1 U3332 ( .A(n4318), .ZN(n7526) );
  AOI22_X1 U3333 ( .A1(reg_mem[1748]), .A2(n4314), .B1(n7530), .B2(data_w[4]), 
        .ZN(n4318) );
  INV_X1 U3334 ( .A(n4319), .ZN(n7527) );
  AOI22_X1 U3335 ( .A1(reg_mem[1749]), .A2(n4314), .B1(n7530), .B2(data_w[5]), 
        .ZN(n4319) );
  INV_X1 U3336 ( .A(n4320), .ZN(n7528) );
  AOI22_X1 U3337 ( .A1(reg_mem[1750]), .A2(n4314), .B1(n7530), .B2(data_w[6]), 
        .ZN(n4320) );
  INV_X1 U3338 ( .A(n4321), .ZN(n7529) );
  AOI22_X1 U3339 ( .A1(reg_mem[1751]), .A2(n4314), .B1(n7530), .B2(data_w[7]), 
        .ZN(n4321) );
  INV_X1 U3340 ( .A(n4322), .ZN(n8099) );
  AOI22_X1 U3341 ( .A1(reg_mem[1752]), .A2(n4323), .B1(n8107), .B2(data_w[0]), 
        .ZN(n4322) );
  INV_X1 U3342 ( .A(n4324), .ZN(n8100) );
  AOI22_X1 U3343 ( .A1(reg_mem[1753]), .A2(n4323), .B1(n8107), .B2(data_w[1]), 
        .ZN(n4324) );
  INV_X1 U3344 ( .A(n4325), .ZN(n8101) );
  AOI22_X1 U3345 ( .A1(reg_mem[1754]), .A2(n4323), .B1(n8107), .B2(data_w[2]), 
        .ZN(n4325) );
  INV_X1 U3346 ( .A(n4326), .ZN(n8102) );
  AOI22_X1 U3347 ( .A1(reg_mem[1755]), .A2(n4323), .B1(n8107), .B2(data_w[3]), 
        .ZN(n4326) );
  INV_X1 U3348 ( .A(n4327), .ZN(n8103) );
  AOI22_X1 U3349 ( .A1(reg_mem[1756]), .A2(n4323), .B1(n8107), .B2(data_w[4]), 
        .ZN(n4327) );
  INV_X1 U3350 ( .A(n4328), .ZN(n8104) );
  AOI22_X1 U3351 ( .A1(reg_mem[1757]), .A2(n4323), .B1(n8107), .B2(data_w[5]), 
        .ZN(n4328) );
  INV_X1 U3352 ( .A(n4329), .ZN(n8105) );
  AOI22_X1 U3353 ( .A1(reg_mem[1758]), .A2(n4323), .B1(n8107), .B2(data_w[6]), 
        .ZN(n4329) );
  INV_X1 U3354 ( .A(n4330), .ZN(n8106) );
  AOI22_X1 U3355 ( .A1(reg_mem[1759]), .A2(n4323), .B1(n8107), .B2(data_w[7]), 
        .ZN(n4330) );
  INV_X1 U3356 ( .A(n4331), .ZN(n6802) );
  AOI22_X1 U3357 ( .A1(reg_mem[1760]), .A2(n4332), .B1(n6810), .B2(data_w[0]), 
        .ZN(n4331) );
  INV_X1 U3358 ( .A(n4333), .ZN(n6803) );
  AOI22_X1 U3359 ( .A1(reg_mem[1761]), .A2(n4332), .B1(n6810), .B2(data_w[1]), 
        .ZN(n4333) );
  INV_X1 U3360 ( .A(n4334), .ZN(n6804) );
  AOI22_X1 U3361 ( .A1(reg_mem[1762]), .A2(n4332), .B1(n6810), .B2(data_w[2]), 
        .ZN(n4334) );
  INV_X1 U3362 ( .A(n4335), .ZN(n6805) );
  AOI22_X1 U3363 ( .A1(reg_mem[1763]), .A2(n4332), .B1(n6810), .B2(data_w[3]), 
        .ZN(n4335) );
  INV_X1 U3364 ( .A(n4336), .ZN(n6806) );
  AOI22_X1 U3365 ( .A1(reg_mem[1764]), .A2(n4332), .B1(n6810), .B2(data_w[4]), 
        .ZN(n4336) );
  INV_X1 U3366 ( .A(n4337), .ZN(n6807) );
  AOI22_X1 U3367 ( .A1(reg_mem[1765]), .A2(n4332), .B1(n6810), .B2(data_w[5]), 
        .ZN(n4337) );
  INV_X1 U3368 ( .A(n4338), .ZN(n6808) );
  AOI22_X1 U3369 ( .A1(reg_mem[1766]), .A2(n4332), .B1(n6810), .B2(data_w[6]), 
        .ZN(n4338) );
  INV_X1 U3370 ( .A(n4339), .ZN(n6809) );
  AOI22_X1 U3371 ( .A1(reg_mem[1767]), .A2(n4332), .B1(n6810), .B2(data_w[7]), 
        .ZN(n4339) );
  INV_X1 U3372 ( .A(n4340), .ZN(n8531) );
  AOI22_X1 U3373 ( .A1(reg_mem[1768]), .A2(n4341), .B1(n8539), .B2(data_w[0]), 
        .ZN(n4340) );
  INV_X1 U3374 ( .A(n4342), .ZN(n8532) );
  AOI22_X1 U3375 ( .A1(reg_mem[1769]), .A2(n4341), .B1(n8539), .B2(data_w[1]), 
        .ZN(n4342) );
  INV_X1 U3376 ( .A(n4343), .ZN(n8533) );
  AOI22_X1 U3377 ( .A1(reg_mem[1770]), .A2(n4341), .B1(n8539), .B2(data_w[2]), 
        .ZN(n4343) );
  INV_X1 U3378 ( .A(n4344), .ZN(n8534) );
  AOI22_X1 U3379 ( .A1(reg_mem[1771]), .A2(n4341), .B1(n8539), .B2(data_w[3]), 
        .ZN(n4344) );
  INV_X1 U3380 ( .A(n4345), .ZN(n8535) );
  AOI22_X1 U3381 ( .A1(reg_mem[1772]), .A2(n4341), .B1(n8539), .B2(data_w[4]), 
        .ZN(n4345) );
  INV_X1 U3382 ( .A(n4346), .ZN(n8536) );
  AOI22_X1 U3383 ( .A1(reg_mem[1773]), .A2(n4341), .B1(n8539), .B2(data_w[5]), 
        .ZN(n4346) );
  INV_X1 U3384 ( .A(n4347), .ZN(n8537) );
  AOI22_X1 U3385 ( .A1(reg_mem[1774]), .A2(n4341), .B1(n8539), .B2(data_w[6]), 
        .ZN(n4347) );
  INV_X1 U3386 ( .A(n4348), .ZN(n8538) );
  AOI22_X1 U3387 ( .A1(reg_mem[1775]), .A2(n4341), .B1(n8539), .B2(data_w[7]), 
        .ZN(n4348) );
  INV_X1 U3388 ( .A(n4349), .ZN(n7378) );
  AOI22_X1 U3389 ( .A1(reg_mem[1776]), .A2(n4350), .B1(n7386), .B2(data_w[0]), 
        .ZN(n4349) );
  INV_X1 U3390 ( .A(n4351), .ZN(n7379) );
  AOI22_X1 U3391 ( .A1(reg_mem[1777]), .A2(n4350), .B1(n7386), .B2(data_w[1]), 
        .ZN(n4351) );
  INV_X1 U3392 ( .A(n4352), .ZN(n7380) );
  AOI22_X1 U3393 ( .A1(reg_mem[1778]), .A2(n4350), .B1(n7386), .B2(data_w[2]), 
        .ZN(n4352) );
  INV_X1 U3394 ( .A(n4353), .ZN(n7381) );
  AOI22_X1 U3395 ( .A1(reg_mem[1779]), .A2(n4350), .B1(n7386), .B2(data_w[3]), 
        .ZN(n4353) );
  INV_X1 U3396 ( .A(n4354), .ZN(n7382) );
  AOI22_X1 U3397 ( .A1(reg_mem[1780]), .A2(n4350), .B1(n7386), .B2(data_w[4]), 
        .ZN(n4354) );
  INV_X1 U3398 ( .A(n4355), .ZN(n7383) );
  AOI22_X1 U3399 ( .A1(reg_mem[1781]), .A2(n4350), .B1(n7386), .B2(data_w[5]), 
        .ZN(n4355) );
  INV_X1 U3400 ( .A(n4356), .ZN(n7384) );
  AOI22_X1 U3401 ( .A1(reg_mem[1782]), .A2(n4350), .B1(n7386), .B2(data_w[6]), 
        .ZN(n4356) );
  INV_X1 U3402 ( .A(n4357), .ZN(n7385) );
  AOI22_X1 U3403 ( .A1(reg_mem[1783]), .A2(n4350), .B1(n7386), .B2(data_w[7]), 
        .ZN(n4357) );
  INV_X1 U3404 ( .A(n4358), .ZN(n7955) );
  AOI22_X1 U3405 ( .A1(reg_mem[1784]), .A2(n4359), .B1(n7963), .B2(data_w[0]), 
        .ZN(n4358) );
  INV_X1 U3406 ( .A(n4360), .ZN(n7956) );
  AOI22_X1 U3407 ( .A1(reg_mem[1785]), .A2(n4359), .B1(n7963), .B2(data_w[1]), 
        .ZN(n4360) );
  INV_X1 U3408 ( .A(n4361), .ZN(n7957) );
  AOI22_X1 U3409 ( .A1(reg_mem[1786]), .A2(n4359), .B1(n7963), .B2(data_w[2]), 
        .ZN(n4361) );
  INV_X1 U3410 ( .A(n4362), .ZN(n7958) );
  AOI22_X1 U3411 ( .A1(reg_mem[1787]), .A2(n4359), .B1(n7963), .B2(data_w[3]), 
        .ZN(n4362) );
  INV_X1 U3412 ( .A(n4363), .ZN(n7959) );
  AOI22_X1 U3413 ( .A1(reg_mem[1788]), .A2(n4359), .B1(n7963), .B2(data_w[4]), 
        .ZN(n4363) );
  INV_X1 U3414 ( .A(n4364), .ZN(n7960) );
  AOI22_X1 U3415 ( .A1(reg_mem[1789]), .A2(n4359), .B1(n7963), .B2(data_w[5]), 
        .ZN(n4364) );
  INV_X1 U3416 ( .A(n4365), .ZN(n7961) );
  AOI22_X1 U3417 ( .A1(reg_mem[1790]), .A2(n4359), .B1(n7963), .B2(data_w[6]), 
        .ZN(n4365) );
  INV_X1 U3418 ( .A(n4366), .ZN(n7962) );
  AOI22_X1 U3419 ( .A1(reg_mem[1791]), .A2(n4359), .B1(n7963), .B2(data_w[7]), 
        .ZN(n4366) );
  INV_X1 U3420 ( .A(n4367), .ZN(n7225) );
  AOI22_X1 U3421 ( .A1(reg_mem[1792]), .A2(n4368), .B1(n7233), .B2(data_w[0]), 
        .ZN(n4367) );
  INV_X1 U3422 ( .A(n4369), .ZN(n7226) );
  AOI22_X1 U3423 ( .A1(reg_mem[1793]), .A2(n4368), .B1(n7233), .B2(data_w[1]), 
        .ZN(n4369) );
  INV_X1 U3424 ( .A(n4370), .ZN(n7227) );
  AOI22_X1 U3425 ( .A1(reg_mem[1794]), .A2(n4368), .B1(n7233), .B2(data_w[2]), 
        .ZN(n4370) );
  INV_X1 U3426 ( .A(n4371), .ZN(n7228) );
  AOI22_X1 U3427 ( .A1(reg_mem[1795]), .A2(n4368), .B1(n7233), .B2(data_w[3]), 
        .ZN(n4371) );
  INV_X1 U3428 ( .A(n4372), .ZN(n7229) );
  AOI22_X1 U3429 ( .A1(reg_mem[1796]), .A2(n4368), .B1(n7233), .B2(data_w[4]), 
        .ZN(n4372) );
  INV_X1 U3430 ( .A(n4373), .ZN(n7230) );
  AOI22_X1 U3431 ( .A1(reg_mem[1797]), .A2(n4368), .B1(n7233), .B2(data_w[5]), 
        .ZN(n4373) );
  INV_X1 U3432 ( .A(n4374), .ZN(n7231) );
  AOI22_X1 U3433 ( .A1(reg_mem[1798]), .A2(n4368), .B1(n7233), .B2(data_w[6]), 
        .ZN(n4374) );
  INV_X1 U3434 ( .A(n4375), .ZN(n7232) );
  AOI22_X1 U3435 ( .A1(reg_mem[1799]), .A2(n4368), .B1(n7233), .B2(data_w[7]), 
        .ZN(n4375) );
  INV_X1 U3436 ( .A(n4377), .ZN(n8954) );
  AOI22_X1 U3437 ( .A1(reg_mem[1800]), .A2(n4378), .B1(n8962), .B2(data_w[0]), 
        .ZN(n4377) );
  INV_X1 U3438 ( .A(n4379), .ZN(n8955) );
  AOI22_X1 U3439 ( .A1(reg_mem[1801]), .A2(n4378), .B1(n8962), .B2(data_w[1]), 
        .ZN(n4379) );
  INV_X1 U3440 ( .A(n4380), .ZN(n8956) );
  AOI22_X1 U3441 ( .A1(reg_mem[1802]), .A2(n4378), .B1(n8962), .B2(data_w[2]), 
        .ZN(n4380) );
  INV_X1 U3442 ( .A(n4381), .ZN(n8957) );
  AOI22_X1 U3443 ( .A1(reg_mem[1803]), .A2(n4378), .B1(n8962), .B2(data_w[3]), 
        .ZN(n4381) );
  INV_X1 U3444 ( .A(n4382), .ZN(n8958) );
  AOI22_X1 U3445 ( .A1(reg_mem[1804]), .A2(n4378), .B1(n8962), .B2(data_w[4]), 
        .ZN(n4382) );
  INV_X1 U3446 ( .A(n4383), .ZN(n8959) );
  AOI22_X1 U3447 ( .A1(reg_mem[1805]), .A2(n4378), .B1(n8962), .B2(data_w[5]), 
        .ZN(n4383) );
  INV_X1 U3448 ( .A(n4384), .ZN(n8960) );
  AOI22_X1 U3449 ( .A1(reg_mem[1806]), .A2(n4378), .B1(n8962), .B2(data_w[6]), 
        .ZN(n4384) );
  INV_X1 U3450 ( .A(n4385), .ZN(n8961) );
  AOI22_X1 U3451 ( .A1(reg_mem[1807]), .A2(n4378), .B1(n8962), .B2(data_w[7]), 
        .ZN(n4385) );
  INV_X1 U3452 ( .A(n4386), .ZN(n7801) );
  AOI22_X1 U3453 ( .A1(reg_mem[1808]), .A2(n4387), .B1(n7809), .B2(data_w[0]), 
        .ZN(n4386) );
  INV_X1 U3454 ( .A(n4388), .ZN(n7802) );
  AOI22_X1 U3455 ( .A1(reg_mem[1809]), .A2(n4387), .B1(n7809), .B2(data_w[1]), 
        .ZN(n4388) );
  INV_X1 U3456 ( .A(n4389), .ZN(n7803) );
  AOI22_X1 U3457 ( .A1(reg_mem[1810]), .A2(n4387), .B1(n7809), .B2(data_w[2]), 
        .ZN(n4389) );
  INV_X1 U3458 ( .A(n4390), .ZN(n7804) );
  AOI22_X1 U3459 ( .A1(reg_mem[1811]), .A2(n4387), .B1(n7809), .B2(data_w[3]), 
        .ZN(n4390) );
  INV_X1 U3460 ( .A(n4391), .ZN(n7805) );
  AOI22_X1 U3461 ( .A1(reg_mem[1812]), .A2(n4387), .B1(n7809), .B2(data_w[4]), 
        .ZN(n4391) );
  INV_X1 U3462 ( .A(n4392), .ZN(n7806) );
  AOI22_X1 U3463 ( .A1(reg_mem[1813]), .A2(n4387), .B1(n7809), .B2(data_w[5]), 
        .ZN(n4392) );
  INV_X1 U3464 ( .A(n4393), .ZN(n7807) );
  AOI22_X1 U3465 ( .A1(reg_mem[1814]), .A2(n4387), .B1(n7809), .B2(data_w[6]), 
        .ZN(n4393) );
  INV_X1 U3466 ( .A(n4394), .ZN(n7808) );
  AOI22_X1 U3467 ( .A1(reg_mem[1815]), .A2(n4387), .B1(n7809), .B2(data_w[7]), 
        .ZN(n4394) );
  INV_X1 U3468 ( .A(n4395), .ZN(n8378) );
  AOI22_X1 U3469 ( .A1(reg_mem[1816]), .A2(n4396), .B1(n8386), .B2(data_w[0]), 
        .ZN(n4395) );
  INV_X1 U3470 ( .A(n4397), .ZN(n8379) );
  AOI22_X1 U3471 ( .A1(reg_mem[1817]), .A2(n4396), .B1(n8386), .B2(data_w[1]), 
        .ZN(n4397) );
  INV_X1 U3472 ( .A(n4398), .ZN(n8380) );
  AOI22_X1 U3473 ( .A1(reg_mem[1818]), .A2(n4396), .B1(n8386), .B2(data_w[2]), 
        .ZN(n4398) );
  INV_X1 U3474 ( .A(n4399), .ZN(n8381) );
  AOI22_X1 U3475 ( .A1(reg_mem[1819]), .A2(n4396), .B1(n8386), .B2(data_w[3]), 
        .ZN(n4399) );
  INV_X1 U3476 ( .A(n4400), .ZN(n8382) );
  AOI22_X1 U3477 ( .A1(reg_mem[1820]), .A2(n4396), .B1(n8386), .B2(data_w[4]), 
        .ZN(n4400) );
  INV_X1 U3478 ( .A(n4401), .ZN(n8383) );
  AOI22_X1 U3479 ( .A1(reg_mem[1821]), .A2(n4396), .B1(n8386), .B2(data_w[5]), 
        .ZN(n4401) );
  INV_X1 U3480 ( .A(n4402), .ZN(n8384) );
  AOI22_X1 U3481 ( .A1(reg_mem[1822]), .A2(n4396), .B1(n8386), .B2(data_w[6]), 
        .ZN(n4402) );
  INV_X1 U3482 ( .A(n4403), .ZN(n8385) );
  AOI22_X1 U3483 ( .A1(reg_mem[1823]), .A2(n4396), .B1(n8386), .B2(data_w[7]), 
        .ZN(n4403) );
  INV_X1 U3484 ( .A(n4404), .ZN(n7081) );
  AOI22_X1 U3485 ( .A1(reg_mem[1824]), .A2(n4405), .B1(n7089), .B2(data_w[0]), 
        .ZN(n4404) );
  INV_X1 U3486 ( .A(n4406), .ZN(n7082) );
  AOI22_X1 U3487 ( .A1(reg_mem[1825]), .A2(n4405), .B1(n7089), .B2(data_w[1]), 
        .ZN(n4406) );
  INV_X1 U3488 ( .A(n4407), .ZN(n7083) );
  AOI22_X1 U3489 ( .A1(reg_mem[1826]), .A2(n4405), .B1(n7089), .B2(data_w[2]), 
        .ZN(n4407) );
  INV_X1 U3490 ( .A(n4408), .ZN(n7084) );
  AOI22_X1 U3491 ( .A1(reg_mem[1827]), .A2(n4405), .B1(n7089), .B2(data_w[3]), 
        .ZN(n4408) );
  INV_X1 U3492 ( .A(n4409), .ZN(n7085) );
  AOI22_X1 U3493 ( .A1(reg_mem[1828]), .A2(n4405), .B1(n7089), .B2(data_w[4]), 
        .ZN(n4409) );
  INV_X1 U3494 ( .A(n4410), .ZN(n7086) );
  AOI22_X1 U3495 ( .A1(reg_mem[1829]), .A2(n4405), .B1(n7089), .B2(data_w[5]), 
        .ZN(n4410) );
  INV_X1 U3496 ( .A(n4411), .ZN(n7087) );
  AOI22_X1 U3497 ( .A1(reg_mem[1830]), .A2(n4405), .B1(n7089), .B2(data_w[6]), 
        .ZN(n4411) );
  INV_X1 U3498 ( .A(n4412), .ZN(n7088) );
  AOI22_X1 U3499 ( .A1(reg_mem[1831]), .A2(n4405), .B1(n7089), .B2(data_w[7]), 
        .ZN(n4412) );
  INV_X1 U3500 ( .A(n4413), .ZN(n8810) );
  AOI22_X1 U3501 ( .A1(reg_mem[1832]), .A2(n4414), .B1(n8818), .B2(data_w[0]), 
        .ZN(n4413) );
  INV_X1 U3502 ( .A(n4415), .ZN(n8811) );
  AOI22_X1 U3503 ( .A1(reg_mem[1833]), .A2(n4414), .B1(n8818), .B2(data_w[1]), 
        .ZN(n4415) );
  INV_X1 U3504 ( .A(n4416), .ZN(n8812) );
  AOI22_X1 U3505 ( .A1(reg_mem[1834]), .A2(n4414), .B1(n8818), .B2(data_w[2]), 
        .ZN(n4416) );
  INV_X1 U3506 ( .A(n4417), .ZN(n8813) );
  AOI22_X1 U3507 ( .A1(reg_mem[1835]), .A2(n4414), .B1(n8818), .B2(data_w[3]), 
        .ZN(n4417) );
  INV_X1 U3508 ( .A(n4418), .ZN(n8814) );
  AOI22_X1 U3509 ( .A1(reg_mem[1836]), .A2(n4414), .B1(n8818), .B2(data_w[4]), 
        .ZN(n4418) );
  INV_X1 U3510 ( .A(n4419), .ZN(n8815) );
  AOI22_X1 U3511 ( .A1(reg_mem[1837]), .A2(n4414), .B1(n8818), .B2(data_w[5]), 
        .ZN(n4419) );
  INV_X1 U3512 ( .A(n4420), .ZN(n8816) );
  AOI22_X1 U3513 ( .A1(reg_mem[1838]), .A2(n4414), .B1(n8818), .B2(data_w[6]), 
        .ZN(n4420) );
  INV_X1 U3514 ( .A(n4421), .ZN(n8817) );
  AOI22_X1 U3515 ( .A1(reg_mem[1839]), .A2(n4414), .B1(n8818), .B2(data_w[7]), 
        .ZN(n4421) );
  INV_X1 U3516 ( .A(n4422), .ZN(n7657) );
  AOI22_X1 U3517 ( .A1(reg_mem[1840]), .A2(n4423), .B1(n7665), .B2(data_w[0]), 
        .ZN(n4422) );
  INV_X1 U3518 ( .A(n4424), .ZN(n7658) );
  AOI22_X1 U3519 ( .A1(reg_mem[1841]), .A2(n4423), .B1(n7665), .B2(data_w[1]), 
        .ZN(n4424) );
  INV_X1 U3520 ( .A(n4425), .ZN(n7659) );
  AOI22_X1 U3521 ( .A1(reg_mem[1842]), .A2(n4423), .B1(n7665), .B2(data_w[2]), 
        .ZN(n4425) );
  INV_X1 U3522 ( .A(n4426), .ZN(n7660) );
  AOI22_X1 U3523 ( .A1(reg_mem[1843]), .A2(n4423), .B1(n7665), .B2(data_w[3]), 
        .ZN(n4426) );
  INV_X1 U3524 ( .A(n4427), .ZN(n7661) );
  AOI22_X1 U3525 ( .A1(reg_mem[1844]), .A2(n4423), .B1(n7665), .B2(data_w[4]), 
        .ZN(n4427) );
  INV_X1 U3526 ( .A(n4428), .ZN(n7662) );
  AOI22_X1 U3527 ( .A1(reg_mem[1845]), .A2(n4423), .B1(n7665), .B2(data_w[5]), 
        .ZN(n4428) );
  INV_X1 U3528 ( .A(n4429), .ZN(n7663) );
  AOI22_X1 U3529 ( .A1(reg_mem[1846]), .A2(n4423), .B1(n7665), .B2(data_w[6]), 
        .ZN(n4429) );
  INV_X1 U3530 ( .A(n4430), .ZN(n7664) );
  AOI22_X1 U3531 ( .A1(reg_mem[1847]), .A2(n4423), .B1(n7665), .B2(data_w[7]), 
        .ZN(n4430) );
  INV_X1 U3532 ( .A(n4431), .ZN(n8234) );
  AOI22_X1 U3533 ( .A1(reg_mem[1848]), .A2(n4432), .B1(n8242), .B2(data_w[0]), 
        .ZN(n4431) );
  INV_X1 U3534 ( .A(n4433), .ZN(n8235) );
  AOI22_X1 U3535 ( .A1(reg_mem[1849]), .A2(n4432), .B1(n8242), .B2(data_w[1]), 
        .ZN(n4433) );
  INV_X1 U3536 ( .A(n4434), .ZN(n8236) );
  AOI22_X1 U3537 ( .A1(reg_mem[1850]), .A2(n4432), .B1(n8242), .B2(data_w[2]), 
        .ZN(n4434) );
  INV_X1 U3538 ( .A(n4435), .ZN(n8237) );
  AOI22_X1 U3539 ( .A1(reg_mem[1851]), .A2(n4432), .B1(n8242), .B2(data_w[3]), 
        .ZN(n4435) );
  INV_X1 U3540 ( .A(n4436), .ZN(n8238) );
  AOI22_X1 U3541 ( .A1(reg_mem[1852]), .A2(n4432), .B1(n8242), .B2(data_w[4]), 
        .ZN(n4436) );
  INV_X1 U3542 ( .A(n4437), .ZN(n8239) );
  AOI22_X1 U3543 ( .A1(reg_mem[1853]), .A2(n4432), .B1(n8242), .B2(data_w[5]), 
        .ZN(n4437) );
  INV_X1 U3544 ( .A(n4438), .ZN(n8240) );
  AOI22_X1 U3545 ( .A1(reg_mem[1854]), .A2(n4432), .B1(n8242), .B2(data_w[6]), 
        .ZN(n4438) );
  INV_X1 U3546 ( .A(n4439), .ZN(n8241) );
  AOI22_X1 U3547 ( .A1(reg_mem[1855]), .A2(n4432), .B1(n8242), .B2(data_w[7]), 
        .ZN(n4439) );
  INV_X1 U3548 ( .A(n4440), .ZN(n6937) );
  AOI22_X1 U3549 ( .A1(reg_mem[1856]), .A2(n4441), .B1(n6945), .B2(data_w[0]), 
        .ZN(n4440) );
  INV_X1 U3550 ( .A(n4442), .ZN(n6938) );
  AOI22_X1 U3551 ( .A1(reg_mem[1857]), .A2(n4441), .B1(n6945), .B2(data_w[1]), 
        .ZN(n4442) );
  INV_X1 U3552 ( .A(n4443), .ZN(n6939) );
  AOI22_X1 U3553 ( .A1(reg_mem[1858]), .A2(n4441), .B1(n6945), .B2(data_w[2]), 
        .ZN(n4443) );
  INV_X1 U3554 ( .A(n4444), .ZN(n6940) );
  AOI22_X1 U3555 ( .A1(reg_mem[1859]), .A2(n4441), .B1(n6945), .B2(data_w[3]), 
        .ZN(n4444) );
  INV_X1 U3556 ( .A(n4445), .ZN(n6941) );
  AOI22_X1 U3557 ( .A1(reg_mem[1860]), .A2(n4441), .B1(n6945), .B2(data_w[4]), 
        .ZN(n4445) );
  INV_X1 U3558 ( .A(n4446), .ZN(n6942) );
  AOI22_X1 U3559 ( .A1(reg_mem[1861]), .A2(n4441), .B1(n6945), .B2(data_w[5]), 
        .ZN(n4446) );
  INV_X1 U3560 ( .A(n4447), .ZN(n6943) );
  AOI22_X1 U3561 ( .A1(reg_mem[1862]), .A2(n4441), .B1(n6945), .B2(data_w[6]), 
        .ZN(n4447) );
  INV_X1 U3562 ( .A(n4448), .ZN(n6944) );
  AOI22_X1 U3563 ( .A1(reg_mem[1863]), .A2(n4441), .B1(n6945), .B2(data_w[7]), 
        .ZN(n4448) );
  INV_X1 U3564 ( .A(n4449), .ZN(n8666) );
  AOI22_X1 U3565 ( .A1(reg_mem[1864]), .A2(n4450), .B1(n8674), .B2(data_w[0]), 
        .ZN(n4449) );
  INV_X1 U3566 ( .A(n4451), .ZN(n8667) );
  AOI22_X1 U3567 ( .A1(reg_mem[1865]), .A2(n4450), .B1(n8674), .B2(data_w[1]), 
        .ZN(n4451) );
  INV_X1 U3568 ( .A(n4452), .ZN(n8668) );
  AOI22_X1 U3569 ( .A1(reg_mem[1866]), .A2(n4450), .B1(n8674), .B2(data_w[2]), 
        .ZN(n4452) );
  INV_X1 U3570 ( .A(n4453), .ZN(n8669) );
  AOI22_X1 U3571 ( .A1(reg_mem[1867]), .A2(n4450), .B1(n8674), .B2(data_w[3]), 
        .ZN(n4453) );
  INV_X1 U3572 ( .A(n4454), .ZN(n8670) );
  AOI22_X1 U3573 ( .A1(reg_mem[1868]), .A2(n4450), .B1(n8674), .B2(data_w[4]), 
        .ZN(n4454) );
  INV_X1 U3574 ( .A(n4455), .ZN(n8671) );
  AOI22_X1 U3575 ( .A1(reg_mem[1869]), .A2(n4450), .B1(n8674), .B2(data_w[5]), 
        .ZN(n4455) );
  INV_X1 U3576 ( .A(n4456), .ZN(n8672) );
  AOI22_X1 U3577 ( .A1(reg_mem[1870]), .A2(n4450), .B1(n8674), .B2(data_w[6]), 
        .ZN(n4456) );
  INV_X1 U3578 ( .A(n4457), .ZN(n8673) );
  AOI22_X1 U3579 ( .A1(reg_mem[1871]), .A2(n4450), .B1(n8674), .B2(data_w[7]), 
        .ZN(n4457) );
  INV_X1 U3580 ( .A(n4458), .ZN(n7513) );
  AOI22_X1 U3581 ( .A1(reg_mem[1872]), .A2(n4459), .B1(n7521), .B2(data_w[0]), 
        .ZN(n4458) );
  INV_X1 U3582 ( .A(n4460), .ZN(n7514) );
  AOI22_X1 U3583 ( .A1(reg_mem[1873]), .A2(n4459), .B1(n7521), .B2(data_w[1]), 
        .ZN(n4460) );
  INV_X1 U3584 ( .A(n4461), .ZN(n7515) );
  AOI22_X1 U3585 ( .A1(reg_mem[1874]), .A2(n4459), .B1(n7521), .B2(data_w[2]), 
        .ZN(n4461) );
  INV_X1 U3586 ( .A(n4462), .ZN(n7516) );
  AOI22_X1 U3587 ( .A1(reg_mem[1875]), .A2(n4459), .B1(n7521), .B2(data_w[3]), 
        .ZN(n4462) );
  INV_X1 U3588 ( .A(n4463), .ZN(n7517) );
  AOI22_X1 U3589 ( .A1(reg_mem[1876]), .A2(n4459), .B1(n7521), .B2(data_w[4]), 
        .ZN(n4463) );
  INV_X1 U3590 ( .A(n4464), .ZN(n7518) );
  AOI22_X1 U3591 ( .A1(reg_mem[1877]), .A2(n4459), .B1(n7521), .B2(data_w[5]), 
        .ZN(n4464) );
  INV_X1 U3592 ( .A(n4465), .ZN(n7519) );
  AOI22_X1 U3593 ( .A1(reg_mem[1878]), .A2(n4459), .B1(n7521), .B2(data_w[6]), 
        .ZN(n4465) );
  INV_X1 U3594 ( .A(n4466), .ZN(n7520) );
  AOI22_X1 U3595 ( .A1(reg_mem[1879]), .A2(n4459), .B1(n7521), .B2(data_w[7]), 
        .ZN(n4466) );
  INV_X1 U3596 ( .A(n4467), .ZN(n8090) );
  AOI22_X1 U3597 ( .A1(reg_mem[1880]), .A2(n4468), .B1(n8098), .B2(data_w[0]), 
        .ZN(n4467) );
  INV_X1 U3598 ( .A(n4469), .ZN(n8091) );
  AOI22_X1 U3599 ( .A1(reg_mem[1881]), .A2(n4468), .B1(n8098), .B2(data_w[1]), 
        .ZN(n4469) );
  INV_X1 U3600 ( .A(n4470), .ZN(n8092) );
  AOI22_X1 U3601 ( .A1(reg_mem[1882]), .A2(n4468), .B1(n8098), .B2(data_w[2]), 
        .ZN(n4470) );
  INV_X1 U3602 ( .A(n4471), .ZN(n8093) );
  AOI22_X1 U3603 ( .A1(reg_mem[1883]), .A2(n4468), .B1(n8098), .B2(data_w[3]), 
        .ZN(n4471) );
  INV_X1 U3604 ( .A(n4472), .ZN(n8094) );
  AOI22_X1 U3605 ( .A1(reg_mem[1884]), .A2(n4468), .B1(n8098), .B2(data_w[4]), 
        .ZN(n4472) );
  INV_X1 U3606 ( .A(n4473), .ZN(n8095) );
  AOI22_X1 U3607 ( .A1(reg_mem[1885]), .A2(n4468), .B1(n8098), .B2(data_w[5]), 
        .ZN(n4473) );
  INV_X1 U3608 ( .A(n4474), .ZN(n8096) );
  AOI22_X1 U3609 ( .A1(reg_mem[1886]), .A2(n4468), .B1(n8098), .B2(data_w[6]), 
        .ZN(n4474) );
  INV_X1 U3610 ( .A(n4475), .ZN(n8097) );
  AOI22_X1 U3611 ( .A1(reg_mem[1887]), .A2(n4468), .B1(n8098), .B2(data_w[7]), 
        .ZN(n4475) );
  INV_X1 U3612 ( .A(n4476), .ZN(n6793) );
  AOI22_X1 U3613 ( .A1(reg_mem[1888]), .A2(n4477), .B1(n6801), .B2(data_w[0]), 
        .ZN(n4476) );
  INV_X1 U3614 ( .A(n4478), .ZN(n6794) );
  AOI22_X1 U3615 ( .A1(reg_mem[1889]), .A2(n4477), .B1(n6801), .B2(data_w[1]), 
        .ZN(n4478) );
  INV_X1 U3616 ( .A(n4479), .ZN(n6795) );
  AOI22_X1 U3617 ( .A1(reg_mem[1890]), .A2(n4477), .B1(n6801), .B2(data_w[2]), 
        .ZN(n4479) );
  INV_X1 U3618 ( .A(n4480), .ZN(n6796) );
  AOI22_X1 U3619 ( .A1(reg_mem[1891]), .A2(n4477), .B1(n6801), .B2(data_w[3]), 
        .ZN(n4480) );
  INV_X1 U3620 ( .A(n4481), .ZN(n6797) );
  AOI22_X1 U3621 ( .A1(reg_mem[1892]), .A2(n4477), .B1(n6801), .B2(data_w[4]), 
        .ZN(n4481) );
  INV_X1 U3622 ( .A(n4482), .ZN(n6798) );
  AOI22_X1 U3623 ( .A1(reg_mem[1893]), .A2(n4477), .B1(n6801), .B2(data_w[5]), 
        .ZN(n4482) );
  INV_X1 U3624 ( .A(n4483), .ZN(n6799) );
  AOI22_X1 U3625 ( .A1(reg_mem[1894]), .A2(n4477), .B1(n6801), .B2(data_w[6]), 
        .ZN(n4483) );
  INV_X1 U3626 ( .A(n4484), .ZN(n6800) );
  AOI22_X1 U3627 ( .A1(reg_mem[1895]), .A2(n4477), .B1(n6801), .B2(data_w[7]), 
        .ZN(n4484) );
  INV_X1 U3628 ( .A(n4485), .ZN(n8522) );
  AOI22_X1 U3629 ( .A1(reg_mem[1896]), .A2(n4486), .B1(n8530), .B2(data_w[0]), 
        .ZN(n4485) );
  INV_X1 U3630 ( .A(n4487), .ZN(n8523) );
  AOI22_X1 U3631 ( .A1(reg_mem[1897]), .A2(n4486), .B1(n8530), .B2(data_w[1]), 
        .ZN(n4487) );
  INV_X1 U3632 ( .A(n4488), .ZN(n8524) );
  AOI22_X1 U3633 ( .A1(reg_mem[1898]), .A2(n4486), .B1(n8530), .B2(data_w[2]), 
        .ZN(n4488) );
  INV_X1 U3634 ( .A(n4489), .ZN(n8525) );
  AOI22_X1 U3635 ( .A1(reg_mem[1899]), .A2(n4486), .B1(n8530), .B2(data_w[3]), 
        .ZN(n4489) );
  INV_X1 U3636 ( .A(n4490), .ZN(n8526) );
  AOI22_X1 U3637 ( .A1(reg_mem[1900]), .A2(n4486), .B1(n8530), .B2(data_w[4]), 
        .ZN(n4490) );
  INV_X1 U3638 ( .A(n4491), .ZN(n8527) );
  AOI22_X1 U3639 ( .A1(reg_mem[1901]), .A2(n4486), .B1(n8530), .B2(data_w[5]), 
        .ZN(n4491) );
  INV_X1 U3640 ( .A(n4492), .ZN(n8528) );
  AOI22_X1 U3641 ( .A1(reg_mem[1902]), .A2(n4486), .B1(n8530), .B2(data_w[6]), 
        .ZN(n4492) );
  INV_X1 U3642 ( .A(n4493), .ZN(n8529) );
  AOI22_X1 U3643 ( .A1(reg_mem[1903]), .A2(n4486), .B1(n8530), .B2(data_w[7]), 
        .ZN(n4493) );
  INV_X1 U3644 ( .A(n4494), .ZN(n7369) );
  AOI22_X1 U3645 ( .A1(reg_mem[1904]), .A2(n4495), .B1(n7377), .B2(data_w[0]), 
        .ZN(n4494) );
  INV_X1 U3646 ( .A(n4496), .ZN(n7370) );
  AOI22_X1 U3647 ( .A1(reg_mem[1905]), .A2(n4495), .B1(n7377), .B2(data_w[1]), 
        .ZN(n4496) );
  INV_X1 U3648 ( .A(n4497), .ZN(n7371) );
  AOI22_X1 U3649 ( .A1(reg_mem[1906]), .A2(n4495), .B1(n7377), .B2(data_w[2]), 
        .ZN(n4497) );
  INV_X1 U3650 ( .A(n4498), .ZN(n7372) );
  AOI22_X1 U3651 ( .A1(reg_mem[1907]), .A2(n4495), .B1(n7377), .B2(data_w[3]), 
        .ZN(n4498) );
  INV_X1 U3652 ( .A(n4499), .ZN(n7373) );
  AOI22_X1 U3653 ( .A1(reg_mem[1908]), .A2(n4495), .B1(n7377), .B2(data_w[4]), 
        .ZN(n4499) );
  INV_X1 U3654 ( .A(n4500), .ZN(n7374) );
  AOI22_X1 U3655 ( .A1(reg_mem[1909]), .A2(n4495), .B1(n7377), .B2(data_w[5]), 
        .ZN(n4500) );
  INV_X1 U3656 ( .A(n4501), .ZN(n7375) );
  AOI22_X1 U3657 ( .A1(reg_mem[1910]), .A2(n4495), .B1(n7377), .B2(data_w[6]), 
        .ZN(n4501) );
  INV_X1 U3658 ( .A(n4502), .ZN(n7376) );
  AOI22_X1 U3659 ( .A1(reg_mem[1911]), .A2(n4495), .B1(n7377), .B2(data_w[7]), 
        .ZN(n4502) );
  INV_X1 U3660 ( .A(n4503), .ZN(n7946) );
  AOI22_X1 U3661 ( .A1(reg_mem[1912]), .A2(n4504), .B1(n7954), .B2(data_w[0]), 
        .ZN(n4503) );
  INV_X1 U3662 ( .A(n4505), .ZN(n7947) );
  AOI22_X1 U3663 ( .A1(reg_mem[1913]), .A2(n4504), .B1(n7954), .B2(data_w[1]), 
        .ZN(n4505) );
  INV_X1 U3664 ( .A(n4506), .ZN(n7948) );
  AOI22_X1 U3665 ( .A1(reg_mem[1914]), .A2(n4504), .B1(n7954), .B2(data_w[2]), 
        .ZN(n4506) );
  INV_X1 U3666 ( .A(n4507), .ZN(n7949) );
  AOI22_X1 U3667 ( .A1(reg_mem[1915]), .A2(n4504), .B1(n7954), .B2(data_w[3]), 
        .ZN(n4507) );
  INV_X1 U3668 ( .A(n4508), .ZN(n7950) );
  AOI22_X1 U3669 ( .A1(reg_mem[1916]), .A2(n4504), .B1(n7954), .B2(data_w[4]), 
        .ZN(n4508) );
  INV_X1 U3670 ( .A(n4509), .ZN(n7951) );
  AOI22_X1 U3671 ( .A1(reg_mem[1917]), .A2(n4504), .B1(n7954), .B2(data_w[5]), 
        .ZN(n4509) );
  INV_X1 U3672 ( .A(n4510), .ZN(n7952) );
  AOI22_X1 U3673 ( .A1(reg_mem[1918]), .A2(n4504), .B1(n7954), .B2(data_w[6]), 
        .ZN(n4510) );
  INV_X1 U3674 ( .A(n4511), .ZN(n7953) );
  AOI22_X1 U3675 ( .A1(reg_mem[1919]), .A2(n4504), .B1(n7954), .B2(data_w[7]), 
        .ZN(n4511) );
  INV_X1 U3676 ( .A(n4512), .ZN(n7216) );
  AOI22_X1 U3677 ( .A1(reg_mem[1920]), .A2(n4513), .B1(n7224), .B2(data_w[0]), 
        .ZN(n4512) );
  INV_X1 U3678 ( .A(n4514), .ZN(n7217) );
  AOI22_X1 U3679 ( .A1(reg_mem[1921]), .A2(n4513), .B1(n7224), .B2(data_w[1]), 
        .ZN(n4514) );
  INV_X1 U3680 ( .A(n4515), .ZN(n7218) );
  AOI22_X1 U3681 ( .A1(reg_mem[1922]), .A2(n4513), .B1(n7224), .B2(data_w[2]), 
        .ZN(n4515) );
  INV_X1 U3682 ( .A(n4516), .ZN(n7219) );
  AOI22_X1 U3683 ( .A1(reg_mem[1923]), .A2(n4513), .B1(n7224), .B2(data_w[3]), 
        .ZN(n4516) );
  INV_X1 U3684 ( .A(n4517), .ZN(n7220) );
  AOI22_X1 U3685 ( .A1(reg_mem[1924]), .A2(n4513), .B1(n7224), .B2(data_w[4]), 
        .ZN(n4517) );
  INV_X1 U3686 ( .A(n4518), .ZN(n7221) );
  AOI22_X1 U3687 ( .A1(reg_mem[1925]), .A2(n4513), .B1(n7224), .B2(data_w[5]), 
        .ZN(n4518) );
  INV_X1 U3688 ( .A(n4519), .ZN(n7222) );
  AOI22_X1 U3689 ( .A1(reg_mem[1926]), .A2(n4513), .B1(n7224), .B2(data_w[6]), 
        .ZN(n4519) );
  INV_X1 U3690 ( .A(n4520), .ZN(n7223) );
  AOI22_X1 U3691 ( .A1(reg_mem[1927]), .A2(n4513), .B1(n7224), .B2(data_w[7]), 
        .ZN(n4520) );
  INV_X1 U3692 ( .A(n4524), .ZN(n8945) );
  AOI22_X1 U3693 ( .A1(reg_mem[1928]), .A2(n4525), .B1(n8953), .B2(data_w[0]), 
        .ZN(n4524) );
  INV_X1 U3694 ( .A(n4526), .ZN(n8946) );
  AOI22_X1 U3695 ( .A1(reg_mem[1929]), .A2(n4525), .B1(n8953), .B2(data_w[1]), 
        .ZN(n4526) );
  INV_X1 U3696 ( .A(n4527), .ZN(n8947) );
  AOI22_X1 U3697 ( .A1(reg_mem[1930]), .A2(n4525), .B1(n8953), .B2(data_w[2]), 
        .ZN(n4527) );
  INV_X1 U3698 ( .A(n4528), .ZN(n8948) );
  AOI22_X1 U3699 ( .A1(reg_mem[1931]), .A2(n4525), .B1(n8953), .B2(data_w[3]), 
        .ZN(n4528) );
  INV_X1 U3700 ( .A(n4529), .ZN(n8949) );
  AOI22_X1 U3701 ( .A1(reg_mem[1932]), .A2(n4525), .B1(n8953), .B2(data_w[4]), 
        .ZN(n4529) );
  INV_X1 U3702 ( .A(n4530), .ZN(n8950) );
  AOI22_X1 U3703 ( .A1(reg_mem[1933]), .A2(n4525), .B1(n8953), .B2(data_w[5]), 
        .ZN(n4530) );
  INV_X1 U3704 ( .A(n4531), .ZN(n8951) );
  AOI22_X1 U3705 ( .A1(reg_mem[1934]), .A2(n4525), .B1(n8953), .B2(data_w[6]), 
        .ZN(n4531) );
  INV_X1 U3706 ( .A(n4532), .ZN(n8952) );
  AOI22_X1 U3707 ( .A1(reg_mem[1935]), .A2(n4525), .B1(n8953), .B2(data_w[7]), 
        .ZN(n4532) );
  INV_X1 U3708 ( .A(n4534), .ZN(n7792) );
  AOI22_X1 U3709 ( .A1(reg_mem[1936]), .A2(n4535), .B1(n7800), .B2(data_w[0]), 
        .ZN(n4534) );
  INV_X1 U3710 ( .A(n4536), .ZN(n7793) );
  AOI22_X1 U3711 ( .A1(reg_mem[1937]), .A2(n4535), .B1(n7800), .B2(data_w[1]), 
        .ZN(n4536) );
  INV_X1 U3712 ( .A(n4537), .ZN(n7794) );
  AOI22_X1 U3713 ( .A1(reg_mem[1938]), .A2(n4535), .B1(n7800), .B2(data_w[2]), 
        .ZN(n4537) );
  INV_X1 U3714 ( .A(n4538), .ZN(n7795) );
  AOI22_X1 U3715 ( .A1(reg_mem[1939]), .A2(n4535), .B1(n7800), .B2(data_w[3]), 
        .ZN(n4538) );
  INV_X1 U3716 ( .A(n4539), .ZN(n7796) );
  AOI22_X1 U3717 ( .A1(reg_mem[1940]), .A2(n4535), .B1(n7800), .B2(data_w[4]), 
        .ZN(n4539) );
  INV_X1 U3718 ( .A(n4540), .ZN(n7797) );
  AOI22_X1 U3719 ( .A1(reg_mem[1941]), .A2(n4535), .B1(n7800), .B2(data_w[5]), 
        .ZN(n4540) );
  INV_X1 U3720 ( .A(n4541), .ZN(n7798) );
  AOI22_X1 U3721 ( .A1(reg_mem[1942]), .A2(n4535), .B1(n7800), .B2(data_w[6]), 
        .ZN(n4541) );
  INV_X1 U3722 ( .A(n4542), .ZN(n7799) );
  AOI22_X1 U3723 ( .A1(reg_mem[1943]), .A2(n4535), .B1(n7800), .B2(data_w[7]), 
        .ZN(n4542) );
  INV_X1 U3724 ( .A(n4544), .ZN(n8369) );
  AOI22_X1 U3725 ( .A1(reg_mem[1944]), .A2(n4545), .B1(n8377), .B2(data_w[0]), 
        .ZN(n4544) );
  INV_X1 U3726 ( .A(n4546), .ZN(n8370) );
  AOI22_X1 U3727 ( .A1(reg_mem[1945]), .A2(n4545), .B1(n8377), .B2(data_w[1]), 
        .ZN(n4546) );
  INV_X1 U3728 ( .A(n4547), .ZN(n8371) );
  AOI22_X1 U3729 ( .A1(reg_mem[1946]), .A2(n4545), .B1(n8377), .B2(data_w[2]), 
        .ZN(n4547) );
  INV_X1 U3730 ( .A(n4548), .ZN(n8372) );
  AOI22_X1 U3731 ( .A1(reg_mem[1947]), .A2(n4545), .B1(n8377), .B2(data_w[3]), 
        .ZN(n4548) );
  INV_X1 U3732 ( .A(n4549), .ZN(n8373) );
  AOI22_X1 U3733 ( .A1(reg_mem[1948]), .A2(n4545), .B1(n8377), .B2(data_w[4]), 
        .ZN(n4549) );
  INV_X1 U3734 ( .A(n4550), .ZN(n8374) );
  AOI22_X1 U3735 ( .A1(reg_mem[1949]), .A2(n4545), .B1(n8377), .B2(data_w[5]), 
        .ZN(n4550) );
  INV_X1 U3736 ( .A(n4551), .ZN(n8375) );
  AOI22_X1 U3737 ( .A1(reg_mem[1950]), .A2(n4545), .B1(n8377), .B2(data_w[6]), 
        .ZN(n4551) );
  INV_X1 U3738 ( .A(n4552), .ZN(n8376) );
  AOI22_X1 U3739 ( .A1(reg_mem[1951]), .A2(n4545), .B1(n8377), .B2(data_w[7]), 
        .ZN(n4552) );
  INV_X1 U3740 ( .A(n4554), .ZN(n7072) );
  AOI22_X1 U3741 ( .A1(reg_mem[1952]), .A2(n4555), .B1(n7080), .B2(data_w[0]), 
        .ZN(n4554) );
  INV_X1 U3742 ( .A(n4556), .ZN(n7073) );
  AOI22_X1 U3743 ( .A1(reg_mem[1953]), .A2(n4555), .B1(n7080), .B2(data_w[1]), 
        .ZN(n4556) );
  INV_X1 U3744 ( .A(n4557), .ZN(n7074) );
  AOI22_X1 U3745 ( .A1(reg_mem[1954]), .A2(n4555), .B1(n7080), .B2(data_w[2]), 
        .ZN(n4557) );
  INV_X1 U3746 ( .A(n4558), .ZN(n7075) );
  AOI22_X1 U3747 ( .A1(reg_mem[1955]), .A2(n4555), .B1(n7080), .B2(data_w[3]), 
        .ZN(n4558) );
  INV_X1 U3748 ( .A(n4559), .ZN(n7076) );
  AOI22_X1 U3749 ( .A1(reg_mem[1956]), .A2(n4555), .B1(n7080), .B2(data_w[4]), 
        .ZN(n4559) );
  INV_X1 U3750 ( .A(n4560), .ZN(n7077) );
  AOI22_X1 U3751 ( .A1(reg_mem[1957]), .A2(n4555), .B1(n7080), .B2(data_w[5]), 
        .ZN(n4560) );
  INV_X1 U3752 ( .A(n4561), .ZN(n7078) );
  AOI22_X1 U3753 ( .A1(reg_mem[1958]), .A2(n4555), .B1(n7080), .B2(data_w[6]), 
        .ZN(n4561) );
  INV_X1 U3754 ( .A(n4562), .ZN(n7079) );
  AOI22_X1 U3755 ( .A1(reg_mem[1959]), .A2(n4555), .B1(n7080), .B2(data_w[7]), 
        .ZN(n4562) );
  INV_X1 U3756 ( .A(n4564), .ZN(n8801) );
  AOI22_X1 U3757 ( .A1(reg_mem[1960]), .A2(n4565), .B1(n8809), .B2(data_w[0]), 
        .ZN(n4564) );
  INV_X1 U3758 ( .A(n4566), .ZN(n8802) );
  AOI22_X1 U3759 ( .A1(reg_mem[1961]), .A2(n4565), .B1(n8809), .B2(data_w[1]), 
        .ZN(n4566) );
  INV_X1 U3760 ( .A(n4567), .ZN(n8803) );
  AOI22_X1 U3761 ( .A1(reg_mem[1962]), .A2(n4565), .B1(n8809), .B2(data_w[2]), 
        .ZN(n4567) );
  INV_X1 U3762 ( .A(n4568), .ZN(n8804) );
  AOI22_X1 U3763 ( .A1(reg_mem[1963]), .A2(n4565), .B1(n8809), .B2(data_w[3]), 
        .ZN(n4568) );
  INV_X1 U3764 ( .A(n4569), .ZN(n8805) );
  AOI22_X1 U3765 ( .A1(reg_mem[1964]), .A2(n4565), .B1(n8809), .B2(data_w[4]), 
        .ZN(n4569) );
  INV_X1 U3766 ( .A(n4570), .ZN(n8806) );
  AOI22_X1 U3767 ( .A1(reg_mem[1965]), .A2(n4565), .B1(n8809), .B2(data_w[5]), 
        .ZN(n4570) );
  INV_X1 U3768 ( .A(n4571), .ZN(n8807) );
  AOI22_X1 U3769 ( .A1(reg_mem[1966]), .A2(n4565), .B1(n8809), .B2(data_w[6]), 
        .ZN(n4571) );
  INV_X1 U3770 ( .A(n4572), .ZN(n8808) );
  AOI22_X1 U3771 ( .A1(reg_mem[1967]), .A2(n4565), .B1(n8809), .B2(data_w[7]), 
        .ZN(n4572) );
  INV_X1 U3772 ( .A(n4573), .ZN(n7648) );
  AOI22_X1 U3773 ( .A1(reg_mem[1968]), .A2(n4574), .B1(n7656), .B2(data_w[0]), 
        .ZN(n4573) );
  INV_X1 U3774 ( .A(n4575), .ZN(n7649) );
  AOI22_X1 U3775 ( .A1(reg_mem[1969]), .A2(n4574), .B1(n7656), .B2(data_w[1]), 
        .ZN(n4575) );
  INV_X1 U3776 ( .A(n4576), .ZN(n7650) );
  AOI22_X1 U3777 ( .A1(reg_mem[1970]), .A2(n4574), .B1(n7656), .B2(data_w[2]), 
        .ZN(n4576) );
  INV_X1 U3778 ( .A(n4577), .ZN(n7651) );
  AOI22_X1 U3779 ( .A1(reg_mem[1971]), .A2(n4574), .B1(n7656), .B2(data_w[3]), 
        .ZN(n4577) );
  INV_X1 U3780 ( .A(n4578), .ZN(n7652) );
  AOI22_X1 U3781 ( .A1(reg_mem[1972]), .A2(n4574), .B1(n7656), .B2(data_w[4]), 
        .ZN(n4578) );
  INV_X1 U3782 ( .A(n4579), .ZN(n7653) );
  AOI22_X1 U3783 ( .A1(reg_mem[1973]), .A2(n4574), .B1(n7656), .B2(data_w[5]), 
        .ZN(n4579) );
  INV_X1 U3784 ( .A(n4580), .ZN(n7654) );
  AOI22_X1 U3785 ( .A1(reg_mem[1974]), .A2(n4574), .B1(n7656), .B2(data_w[6]), 
        .ZN(n4580) );
  INV_X1 U3786 ( .A(n4581), .ZN(n7655) );
  AOI22_X1 U3787 ( .A1(reg_mem[1975]), .A2(n4574), .B1(n7656), .B2(data_w[7]), 
        .ZN(n4581) );
  INV_X1 U3788 ( .A(n4582), .ZN(n8225) );
  AOI22_X1 U3789 ( .A1(reg_mem[1976]), .A2(n4583), .B1(n8233), .B2(data_w[0]), 
        .ZN(n4582) );
  INV_X1 U3790 ( .A(n4584), .ZN(n8226) );
  AOI22_X1 U3791 ( .A1(reg_mem[1977]), .A2(n4583), .B1(n8233), .B2(data_w[1]), 
        .ZN(n4584) );
  INV_X1 U3792 ( .A(n4585), .ZN(n8227) );
  AOI22_X1 U3793 ( .A1(reg_mem[1978]), .A2(n4583), .B1(n8233), .B2(data_w[2]), 
        .ZN(n4585) );
  INV_X1 U3794 ( .A(n4586), .ZN(n8228) );
  AOI22_X1 U3795 ( .A1(reg_mem[1979]), .A2(n4583), .B1(n8233), .B2(data_w[3]), 
        .ZN(n4586) );
  INV_X1 U3796 ( .A(n4587), .ZN(n8229) );
  AOI22_X1 U3797 ( .A1(reg_mem[1980]), .A2(n4583), .B1(n8233), .B2(data_w[4]), 
        .ZN(n4587) );
  INV_X1 U3798 ( .A(n4588), .ZN(n8230) );
  AOI22_X1 U3799 ( .A1(reg_mem[1981]), .A2(n4583), .B1(n8233), .B2(data_w[5]), 
        .ZN(n4588) );
  INV_X1 U3800 ( .A(n4589), .ZN(n8231) );
  AOI22_X1 U3801 ( .A1(reg_mem[1982]), .A2(n4583), .B1(n8233), .B2(data_w[6]), 
        .ZN(n4589) );
  INV_X1 U3802 ( .A(n4590), .ZN(n8232) );
  AOI22_X1 U3803 ( .A1(reg_mem[1983]), .A2(n4583), .B1(n8233), .B2(data_w[7]), 
        .ZN(n4590) );
  INV_X1 U3804 ( .A(n4591), .ZN(n6928) );
  AOI22_X1 U3805 ( .A1(reg_mem[1984]), .A2(n4592), .B1(n6936), .B2(data_w[0]), 
        .ZN(n4591) );
  INV_X1 U3806 ( .A(n4593), .ZN(n6929) );
  AOI22_X1 U3807 ( .A1(reg_mem[1985]), .A2(n4592), .B1(n6936), .B2(data_w[1]), 
        .ZN(n4593) );
  INV_X1 U3808 ( .A(n4594), .ZN(n6930) );
  AOI22_X1 U3809 ( .A1(reg_mem[1986]), .A2(n4592), .B1(n6936), .B2(data_w[2]), 
        .ZN(n4594) );
  INV_X1 U3810 ( .A(n4595), .ZN(n6931) );
  AOI22_X1 U3811 ( .A1(reg_mem[1987]), .A2(n4592), .B1(n6936), .B2(data_w[3]), 
        .ZN(n4595) );
  INV_X1 U3812 ( .A(n4596), .ZN(n6932) );
  AOI22_X1 U3813 ( .A1(reg_mem[1988]), .A2(n4592), .B1(n6936), .B2(data_w[4]), 
        .ZN(n4596) );
  INV_X1 U3814 ( .A(n4597), .ZN(n6933) );
  AOI22_X1 U3815 ( .A1(reg_mem[1989]), .A2(n4592), .B1(n6936), .B2(data_w[5]), 
        .ZN(n4597) );
  INV_X1 U3816 ( .A(n4598), .ZN(n6934) );
  AOI22_X1 U3817 ( .A1(reg_mem[1990]), .A2(n4592), .B1(n6936), .B2(data_w[6]), 
        .ZN(n4598) );
  INV_X1 U3818 ( .A(n4599), .ZN(n6935) );
  AOI22_X1 U3819 ( .A1(reg_mem[1991]), .A2(n4592), .B1(n6936), .B2(data_w[7]), 
        .ZN(n4599) );
  INV_X1 U3820 ( .A(n4601), .ZN(n8657) );
  AOI22_X1 U3821 ( .A1(reg_mem[1992]), .A2(n4602), .B1(n8665), .B2(data_w[0]), 
        .ZN(n4601) );
  INV_X1 U3822 ( .A(n4603), .ZN(n8658) );
  AOI22_X1 U3823 ( .A1(reg_mem[1993]), .A2(n4602), .B1(n8665), .B2(data_w[1]), 
        .ZN(n4603) );
  INV_X1 U3824 ( .A(n4604), .ZN(n8659) );
  AOI22_X1 U3825 ( .A1(reg_mem[1994]), .A2(n4602), .B1(n8665), .B2(data_w[2]), 
        .ZN(n4604) );
  INV_X1 U3826 ( .A(n4605), .ZN(n8660) );
  AOI22_X1 U3827 ( .A1(reg_mem[1995]), .A2(n4602), .B1(n8665), .B2(data_w[3]), 
        .ZN(n4605) );
  INV_X1 U3828 ( .A(n4606), .ZN(n8661) );
  AOI22_X1 U3829 ( .A1(reg_mem[1996]), .A2(n4602), .B1(n8665), .B2(data_w[4]), 
        .ZN(n4606) );
  INV_X1 U3830 ( .A(n4607), .ZN(n8662) );
  AOI22_X1 U3831 ( .A1(reg_mem[1997]), .A2(n4602), .B1(n8665), .B2(data_w[5]), 
        .ZN(n4607) );
  INV_X1 U3832 ( .A(n4608), .ZN(n8663) );
  AOI22_X1 U3833 ( .A1(reg_mem[1998]), .A2(n4602), .B1(n8665), .B2(data_w[6]), 
        .ZN(n4608) );
  INV_X1 U3834 ( .A(n4609), .ZN(n8664) );
  AOI22_X1 U3835 ( .A1(reg_mem[1999]), .A2(n4602), .B1(n8665), .B2(data_w[7]), 
        .ZN(n4609) );
  INV_X1 U3836 ( .A(n4610), .ZN(n7504) );
  AOI22_X1 U3837 ( .A1(reg_mem[2000]), .A2(n4611), .B1(n7512), .B2(data_w[0]), 
        .ZN(n4610) );
  INV_X1 U3838 ( .A(n4612), .ZN(n7505) );
  AOI22_X1 U3839 ( .A1(reg_mem[2001]), .A2(n4611), .B1(n7512), .B2(data_w[1]), 
        .ZN(n4612) );
  INV_X1 U3840 ( .A(n4613), .ZN(n7506) );
  AOI22_X1 U3841 ( .A1(reg_mem[2002]), .A2(n4611), .B1(n7512), .B2(data_w[2]), 
        .ZN(n4613) );
  INV_X1 U3842 ( .A(n4614), .ZN(n7507) );
  AOI22_X1 U3843 ( .A1(reg_mem[2003]), .A2(n4611), .B1(n7512), .B2(data_w[3]), 
        .ZN(n4614) );
  INV_X1 U3844 ( .A(n4615), .ZN(n7508) );
  AOI22_X1 U3845 ( .A1(reg_mem[2004]), .A2(n4611), .B1(n7512), .B2(data_w[4]), 
        .ZN(n4615) );
  INV_X1 U3846 ( .A(n4616), .ZN(n7509) );
  AOI22_X1 U3847 ( .A1(reg_mem[2005]), .A2(n4611), .B1(n7512), .B2(data_w[5]), 
        .ZN(n4616) );
  INV_X1 U3848 ( .A(n4617), .ZN(n7510) );
  AOI22_X1 U3849 ( .A1(reg_mem[2006]), .A2(n4611), .B1(n7512), .B2(data_w[6]), 
        .ZN(n4617) );
  INV_X1 U3850 ( .A(n4618), .ZN(n7511) );
  AOI22_X1 U3851 ( .A1(reg_mem[2007]), .A2(n4611), .B1(n7512), .B2(data_w[7]), 
        .ZN(n4618) );
  INV_X1 U3852 ( .A(n4619), .ZN(n8081) );
  AOI22_X1 U3853 ( .A1(reg_mem[2008]), .A2(n4620), .B1(n8089), .B2(data_w[0]), 
        .ZN(n4619) );
  INV_X1 U3854 ( .A(n4621), .ZN(n8082) );
  AOI22_X1 U3855 ( .A1(reg_mem[2009]), .A2(n4620), .B1(n8089), .B2(data_w[1]), 
        .ZN(n4621) );
  INV_X1 U3856 ( .A(n4622), .ZN(n8083) );
  AOI22_X1 U3857 ( .A1(reg_mem[2010]), .A2(n4620), .B1(n8089), .B2(data_w[2]), 
        .ZN(n4622) );
  INV_X1 U3858 ( .A(n4623), .ZN(n8084) );
  AOI22_X1 U3859 ( .A1(reg_mem[2011]), .A2(n4620), .B1(n8089), .B2(data_w[3]), 
        .ZN(n4623) );
  INV_X1 U3860 ( .A(n4624), .ZN(n8085) );
  AOI22_X1 U3861 ( .A1(reg_mem[2012]), .A2(n4620), .B1(n8089), .B2(data_w[4]), 
        .ZN(n4624) );
  INV_X1 U3862 ( .A(n4625), .ZN(n8086) );
  AOI22_X1 U3863 ( .A1(reg_mem[2013]), .A2(n4620), .B1(n8089), .B2(data_w[5]), 
        .ZN(n4625) );
  INV_X1 U3864 ( .A(n4626), .ZN(n8087) );
  AOI22_X1 U3865 ( .A1(reg_mem[2014]), .A2(n4620), .B1(n8089), .B2(data_w[6]), 
        .ZN(n4626) );
  INV_X1 U3866 ( .A(n4627), .ZN(n8088) );
  AOI22_X1 U3867 ( .A1(reg_mem[2015]), .A2(n4620), .B1(n8089), .B2(data_w[7]), 
        .ZN(n4627) );
  INV_X1 U3868 ( .A(n4628), .ZN(n6784) );
  AOI22_X1 U3869 ( .A1(reg_mem[2016]), .A2(n4629), .B1(n6792), .B2(data_w[0]), 
        .ZN(n4628) );
  INV_X1 U3870 ( .A(n4630), .ZN(n6785) );
  AOI22_X1 U3871 ( .A1(reg_mem[2017]), .A2(n4629), .B1(n6792), .B2(data_w[1]), 
        .ZN(n4630) );
  INV_X1 U3872 ( .A(n4631), .ZN(n6786) );
  AOI22_X1 U3873 ( .A1(reg_mem[2018]), .A2(n4629), .B1(n6792), .B2(data_w[2]), 
        .ZN(n4631) );
  INV_X1 U3874 ( .A(n4632), .ZN(n6787) );
  AOI22_X1 U3875 ( .A1(reg_mem[2019]), .A2(n4629), .B1(n6792), .B2(data_w[3]), 
        .ZN(n4632) );
  INV_X1 U3876 ( .A(n4633), .ZN(n6788) );
  AOI22_X1 U3877 ( .A1(reg_mem[2020]), .A2(n4629), .B1(n6792), .B2(data_w[4]), 
        .ZN(n4633) );
  INV_X1 U3878 ( .A(n4634), .ZN(n6789) );
  AOI22_X1 U3879 ( .A1(reg_mem[2021]), .A2(n4629), .B1(n6792), .B2(data_w[5]), 
        .ZN(n4634) );
  INV_X1 U3880 ( .A(n4635), .ZN(n6790) );
  AOI22_X1 U3881 ( .A1(reg_mem[2022]), .A2(n4629), .B1(n6792), .B2(data_w[6]), 
        .ZN(n4635) );
  INV_X1 U3882 ( .A(n4636), .ZN(n6791) );
  AOI22_X1 U3883 ( .A1(reg_mem[2023]), .A2(n4629), .B1(n6792), .B2(data_w[7]), 
        .ZN(n4636) );
  INV_X1 U3884 ( .A(n4638), .ZN(n8513) );
  AOI22_X1 U3885 ( .A1(reg_mem[2024]), .A2(n4639), .B1(n8521), .B2(data_w[0]), 
        .ZN(n4638) );
  INV_X1 U3886 ( .A(n4640), .ZN(n8514) );
  AOI22_X1 U3887 ( .A1(reg_mem[2025]), .A2(n4639), .B1(n8521), .B2(data_w[1]), 
        .ZN(n4640) );
  INV_X1 U3888 ( .A(n4641), .ZN(n8515) );
  AOI22_X1 U3889 ( .A1(reg_mem[2026]), .A2(n4639), .B1(n8521), .B2(data_w[2]), 
        .ZN(n4641) );
  INV_X1 U3890 ( .A(n4642), .ZN(n8516) );
  AOI22_X1 U3891 ( .A1(reg_mem[2027]), .A2(n4639), .B1(n8521), .B2(data_w[3]), 
        .ZN(n4642) );
  INV_X1 U3892 ( .A(n4643), .ZN(n8517) );
  AOI22_X1 U3893 ( .A1(reg_mem[2028]), .A2(n4639), .B1(n8521), .B2(data_w[4]), 
        .ZN(n4643) );
  INV_X1 U3894 ( .A(n4644), .ZN(n8518) );
  AOI22_X1 U3895 ( .A1(reg_mem[2029]), .A2(n4639), .B1(n8521), .B2(data_w[5]), 
        .ZN(n4644) );
  INV_X1 U3896 ( .A(n4645), .ZN(n8519) );
  AOI22_X1 U3897 ( .A1(reg_mem[2030]), .A2(n4639), .B1(n8521), .B2(data_w[6]), 
        .ZN(n4645) );
  INV_X1 U3898 ( .A(n4646), .ZN(n8520) );
  AOI22_X1 U3899 ( .A1(reg_mem[2031]), .A2(n4639), .B1(n8521), .B2(data_w[7]), 
        .ZN(n4646) );
  INV_X1 U3900 ( .A(n4647), .ZN(n7360) );
  AOI22_X1 U3901 ( .A1(reg_mem[2032]), .A2(n4648), .B1(n7368), .B2(data_w[0]), 
        .ZN(n4647) );
  INV_X1 U3902 ( .A(n4649), .ZN(n7361) );
  AOI22_X1 U3903 ( .A1(reg_mem[2033]), .A2(n4648), .B1(n7368), .B2(data_w[1]), 
        .ZN(n4649) );
  INV_X1 U3904 ( .A(n4650), .ZN(n7362) );
  AOI22_X1 U3905 ( .A1(reg_mem[2034]), .A2(n4648), .B1(n7368), .B2(data_w[2]), 
        .ZN(n4650) );
  INV_X1 U3906 ( .A(n4651), .ZN(n7363) );
  AOI22_X1 U3907 ( .A1(reg_mem[2035]), .A2(n4648), .B1(n7368), .B2(data_w[3]), 
        .ZN(n4651) );
  INV_X1 U3908 ( .A(n4652), .ZN(n7364) );
  AOI22_X1 U3909 ( .A1(reg_mem[2036]), .A2(n4648), .B1(n7368), .B2(data_w[4]), 
        .ZN(n4652) );
  INV_X1 U3910 ( .A(n4653), .ZN(n7365) );
  AOI22_X1 U3911 ( .A1(reg_mem[2037]), .A2(n4648), .B1(n7368), .B2(data_w[5]), 
        .ZN(n4653) );
  INV_X1 U3912 ( .A(n4654), .ZN(n7366) );
  AOI22_X1 U3913 ( .A1(reg_mem[2038]), .A2(n4648), .B1(n7368), .B2(data_w[6]), 
        .ZN(n4654) );
  INV_X1 U3914 ( .A(n4655), .ZN(n7367) );
  AOI22_X1 U3915 ( .A1(reg_mem[2039]), .A2(n4648), .B1(n7368), .B2(data_w[7]), 
        .ZN(n4655) );
  INV_X1 U3916 ( .A(n4656), .ZN(n7937) );
  AOI22_X1 U3917 ( .A1(reg_mem[2040]), .A2(n4657), .B1(n7945), .B2(data_w[0]), 
        .ZN(n4656) );
  INV_X1 U3918 ( .A(n4658), .ZN(n7938) );
  AOI22_X1 U3919 ( .A1(reg_mem[2041]), .A2(n4657), .B1(n7945), .B2(data_w[1]), 
        .ZN(n4658) );
  INV_X1 U3920 ( .A(n4659), .ZN(n7939) );
  AOI22_X1 U3921 ( .A1(reg_mem[2042]), .A2(n4657), .B1(n7945), .B2(data_w[2]), 
        .ZN(n4659) );
  INV_X1 U3922 ( .A(n4660), .ZN(n7940) );
  AOI22_X1 U3923 ( .A1(reg_mem[2043]), .A2(n4657), .B1(n7945), .B2(data_w[3]), 
        .ZN(n4660) );
  INV_X1 U3924 ( .A(n4661), .ZN(n7941) );
  AOI22_X1 U3925 ( .A1(reg_mem[2044]), .A2(n4657), .B1(n7945), .B2(data_w[4]), 
        .ZN(n4661) );
  INV_X1 U3926 ( .A(n4662), .ZN(n7942) );
  AOI22_X1 U3927 ( .A1(reg_mem[2045]), .A2(n4657), .B1(n7945), .B2(data_w[5]), 
        .ZN(n4662) );
  INV_X1 U3928 ( .A(n4663), .ZN(n7943) );
  AOI22_X1 U3929 ( .A1(reg_mem[2046]), .A2(n4657), .B1(n7945), .B2(data_w[6]), 
        .ZN(n4663) );
  INV_X1 U3930 ( .A(n4664), .ZN(n7944) );
  AOI22_X1 U3931 ( .A1(reg_mem[2047]), .A2(n4657), .B1(n7945), .B2(data_w[7]), 
        .ZN(n4664) );
  INV_X1 U3932 ( .A(n2313), .ZN(n7351) );
  AOI22_X1 U3933 ( .A1(reg_mem[0]), .A2(n2314), .B1(data_w[0]), .B2(n7359), 
        .ZN(n2313) );
  INV_X1 U3934 ( .A(n2315), .ZN(n7352) );
  AOI22_X1 U3935 ( .A1(reg_mem[1]), .A2(n2314), .B1(data_w[1]), .B2(n7359), 
        .ZN(n2315) );
  INV_X1 U3936 ( .A(n2316), .ZN(n7353) );
  AOI22_X1 U3937 ( .A1(reg_mem[2]), .A2(n2314), .B1(data_w[2]), .B2(n7359), 
        .ZN(n2316) );
  INV_X1 U3938 ( .A(n2317), .ZN(n7354) );
  AOI22_X1 U3939 ( .A1(reg_mem[3]), .A2(n2314), .B1(data_w[3]), .B2(n7359), 
        .ZN(n2317) );
  INV_X1 U3940 ( .A(n2318), .ZN(n7355) );
  AOI22_X1 U3941 ( .A1(reg_mem[4]), .A2(n2314), .B1(data_w[4]), .B2(n7359), 
        .ZN(n2318) );
  INV_X1 U3942 ( .A(n2319), .ZN(n7356) );
  AOI22_X1 U3943 ( .A1(reg_mem[5]), .A2(n2314), .B1(data_w[5]), .B2(n7359), 
        .ZN(n2319) );
  INV_X1 U3944 ( .A(n2320), .ZN(n7357) );
  AOI22_X1 U3945 ( .A1(reg_mem[6]), .A2(n2314), .B1(data_w[6]), .B2(n7359), 
        .ZN(n2320) );
  INV_X1 U3946 ( .A(n2321), .ZN(n7358) );
  AOI22_X1 U3947 ( .A1(reg_mem[7]), .A2(n2314), .B1(data_w[7]), .B2(n7359), 
        .ZN(n2321) );
  INV_X1 U3948 ( .A(n2354), .ZN(n7207) );
  AOI22_X1 U3949 ( .A1(reg_mem[32]), .A2(n2355), .B1(n7215), .B2(data_w[0]), 
        .ZN(n2354) );
  INV_X1 U3950 ( .A(n2356), .ZN(n7208) );
  AOI22_X1 U3951 ( .A1(reg_mem[33]), .A2(n2355), .B1(n7215), .B2(data_w[1]), 
        .ZN(n2356) );
  INV_X1 U3952 ( .A(n2357), .ZN(n7209) );
  AOI22_X1 U3953 ( .A1(reg_mem[34]), .A2(n2355), .B1(n7215), .B2(data_w[2]), 
        .ZN(n2357) );
  INV_X1 U3954 ( .A(n2358), .ZN(n7210) );
  AOI22_X1 U3955 ( .A1(reg_mem[35]), .A2(n2355), .B1(n7215), .B2(data_w[3]), 
        .ZN(n2358) );
  INV_X1 U3956 ( .A(n2359), .ZN(n7211) );
  AOI22_X1 U3957 ( .A1(reg_mem[36]), .A2(n2355), .B1(n7215), .B2(data_w[4]), 
        .ZN(n2359) );
  INV_X1 U3958 ( .A(n2360), .ZN(n7212) );
  AOI22_X1 U3959 ( .A1(reg_mem[37]), .A2(n2355), .B1(n7215), .B2(data_w[5]), 
        .ZN(n2360) );
  INV_X1 U3960 ( .A(n2361), .ZN(n7213) );
  AOI22_X1 U3961 ( .A1(reg_mem[38]), .A2(n2355), .B1(n7215), .B2(data_w[6]), 
        .ZN(n2361) );
  INV_X1 U3962 ( .A(n2362), .ZN(n7214) );
  AOI22_X1 U3963 ( .A1(reg_mem[39]), .A2(n2355), .B1(n7215), .B2(data_w[7]), 
        .ZN(n2362) );
  INV_X1 U3964 ( .A(n2364), .ZN(n8936) );
  AOI22_X1 U3965 ( .A1(reg_mem[40]), .A2(n2365), .B1(n8944), .B2(data_w[0]), 
        .ZN(n2364) );
  INV_X1 U3966 ( .A(n2366), .ZN(n8937) );
  AOI22_X1 U3967 ( .A1(reg_mem[41]), .A2(n2365), .B1(n8944), .B2(data_w[1]), 
        .ZN(n2366) );
  INV_X1 U3968 ( .A(n2367), .ZN(n8938) );
  AOI22_X1 U3969 ( .A1(reg_mem[42]), .A2(n2365), .B1(n8944), .B2(data_w[2]), 
        .ZN(n2367) );
  INV_X1 U3970 ( .A(n2368), .ZN(n8939) );
  AOI22_X1 U3971 ( .A1(reg_mem[43]), .A2(n2365), .B1(n8944), .B2(data_w[3]), 
        .ZN(n2368) );
  INV_X1 U3972 ( .A(n2369), .ZN(n8940) );
  AOI22_X1 U3973 ( .A1(reg_mem[44]), .A2(n2365), .B1(n8944), .B2(data_w[4]), 
        .ZN(n2369) );
  INV_X1 U3974 ( .A(n2370), .ZN(n8941) );
  AOI22_X1 U3975 ( .A1(reg_mem[45]), .A2(n2365), .B1(n8944), .B2(data_w[5]), 
        .ZN(n2370) );
  INV_X1 U3976 ( .A(n2371), .ZN(n8942) );
  AOI22_X1 U3977 ( .A1(reg_mem[46]), .A2(n2365), .B1(n8944), .B2(data_w[6]), 
        .ZN(n2371) );
  INV_X1 U3978 ( .A(n2372), .ZN(n8943) );
  AOI22_X1 U3979 ( .A1(reg_mem[47]), .A2(n2365), .B1(n8944), .B2(data_w[7]), 
        .ZN(n2372) );
  INV_X1 U3980 ( .A(n2374), .ZN(n7783) );
  AOI22_X1 U3981 ( .A1(reg_mem[48]), .A2(n2375), .B1(n7791), .B2(data_w[0]), 
        .ZN(n2374) );
  INV_X1 U3982 ( .A(n2376), .ZN(n7784) );
  AOI22_X1 U3983 ( .A1(reg_mem[49]), .A2(n2375), .B1(n7791), .B2(data_w[1]), 
        .ZN(n2376) );
  INV_X1 U3984 ( .A(n2377), .ZN(n7785) );
  AOI22_X1 U3985 ( .A1(reg_mem[50]), .A2(n2375), .B1(n7791), .B2(data_w[2]), 
        .ZN(n2377) );
  INV_X1 U3986 ( .A(n2378), .ZN(n7786) );
  AOI22_X1 U3987 ( .A1(reg_mem[51]), .A2(n2375), .B1(n7791), .B2(data_w[3]), 
        .ZN(n2378) );
  INV_X1 U3988 ( .A(n2379), .ZN(n7787) );
  AOI22_X1 U3989 ( .A1(reg_mem[52]), .A2(n2375), .B1(n7791), .B2(data_w[4]), 
        .ZN(n2379) );
  INV_X1 U3990 ( .A(n2380), .ZN(n7788) );
  AOI22_X1 U3991 ( .A1(reg_mem[53]), .A2(n2375), .B1(n7791), .B2(data_w[5]), 
        .ZN(n2380) );
  INV_X1 U3992 ( .A(n2381), .ZN(n7789) );
  AOI22_X1 U3993 ( .A1(reg_mem[54]), .A2(n2375), .B1(n7791), .B2(data_w[6]), 
        .ZN(n2381) );
  INV_X1 U3994 ( .A(n2382), .ZN(n7790) );
  AOI22_X1 U3995 ( .A1(reg_mem[55]), .A2(n2375), .B1(n7791), .B2(data_w[7]), 
        .ZN(n2382) );
  INV_X1 U3996 ( .A(n2384), .ZN(n8360) );
  AOI22_X1 U3997 ( .A1(reg_mem[56]), .A2(n2385), .B1(n8368), .B2(data_w[0]), 
        .ZN(n2384) );
  INV_X1 U3998 ( .A(n2386), .ZN(n8361) );
  AOI22_X1 U3999 ( .A1(reg_mem[57]), .A2(n2385), .B1(n8368), .B2(data_w[1]), 
        .ZN(n2386) );
  INV_X1 U4000 ( .A(n2387), .ZN(n8362) );
  AOI22_X1 U4001 ( .A1(reg_mem[58]), .A2(n2385), .B1(n8368), .B2(data_w[2]), 
        .ZN(n2387) );
  INV_X1 U4002 ( .A(n2388), .ZN(n8363) );
  AOI22_X1 U4003 ( .A1(reg_mem[59]), .A2(n2385), .B1(n8368), .B2(data_w[3]), 
        .ZN(n2388) );
  INV_X1 U4004 ( .A(n2389), .ZN(n8364) );
  AOI22_X1 U4005 ( .A1(reg_mem[60]), .A2(n2385), .B1(n8368), .B2(data_w[4]), 
        .ZN(n2389) );
  INV_X1 U4006 ( .A(n2390), .ZN(n8365) );
  AOI22_X1 U4007 ( .A1(reg_mem[61]), .A2(n2385), .B1(n8368), .B2(data_w[5]), 
        .ZN(n2390) );
  INV_X1 U4008 ( .A(n2391), .ZN(n8366) );
  AOI22_X1 U4009 ( .A1(reg_mem[62]), .A2(n2385), .B1(n8368), .B2(data_w[6]), 
        .ZN(n2391) );
  INV_X1 U4010 ( .A(n2392), .ZN(n8367) );
  AOI22_X1 U4011 ( .A1(reg_mem[63]), .A2(n2385), .B1(n8368), .B2(data_w[7]), 
        .ZN(n2392) );
  INV_X1 U4012 ( .A(n2394), .ZN(n7063) );
  AOI22_X1 U4013 ( .A1(reg_mem[64]), .A2(n2395), .B1(n7071), .B2(data_w[0]), 
        .ZN(n2394) );
  INV_X1 U4014 ( .A(n2396), .ZN(n7064) );
  AOI22_X1 U4015 ( .A1(reg_mem[65]), .A2(n2395), .B1(n7071), .B2(data_w[1]), 
        .ZN(n2396) );
  INV_X1 U4016 ( .A(n2397), .ZN(n7065) );
  AOI22_X1 U4017 ( .A1(reg_mem[66]), .A2(n2395), .B1(n7071), .B2(data_w[2]), 
        .ZN(n2397) );
  INV_X1 U4018 ( .A(n2398), .ZN(n7066) );
  AOI22_X1 U4019 ( .A1(reg_mem[67]), .A2(n2395), .B1(n7071), .B2(data_w[3]), 
        .ZN(n2398) );
  INV_X1 U4020 ( .A(n2399), .ZN(n7067) );
  AOI22_X1 U4021 ( .A1(reg_mem[68]), .A2(n2395), .B1(n7071), .B2(data_w[4]), 
        .ZN(n2399) );
  INV_X1 U4022 ( .A(n2400), .ZN(n7068) );
  AOI22_X1 U4023 ( .A1(reg_mem[69]), .A2(n2395), .B1(n7071), .B2(data_w[5]), 
        .ZN(n2400) );
  INV_X1 U4024 ( .A(n2401), .ZN(n7069) );
  AOI22_X1 U4025 ( .A1(reg_mem[70]), .A2(n2395), .B1(n7071), .B2(data_w[6]), 
        .ZN(n2401) );
  INV_X1 U4026 ( .A(n2402), .ZN(n7070) );
  AOI22_X1 U4027 ( .A1(reg_mem[71]), .A2(n2395), .B1(n7071), .B2(data_w[7]), 
        .ZN(n2402) );
  INV_X1 U4028 ( .A(n2404), .ZN(n8792) );
  AOI22_X1 U4029 ( .A1(reg_mem[72]), .A2(n2405), .B1(n8800), .B2(data_w[0]), 
        .ZN(n2404) );
  INV_X1 U4030 ( .A(n2406), .ZN(n8793) );
  AOI22_X1 U4031 ( .A1(reg_mem[73]), .A2(n2405), .B1(n8800), .B2(data_w[1]), 
        .ZN(n2406) );
  INV_X1 U4032 ( .A(n2407), .ZN(n8794) );
  AOI22_X1 U4033 ( .A1(reg_mem[74]), .A2(n2405), .B1(n8800), .B2(data_w[2]), 
        .ZN(n2407) );
  INV_X1 U4034 ( .A(n2408), .ZN(n8795) );
  AOI22_X1 U4035 ( .A1(reg_mem[75]), .A2(n2405), .B1(n8800), .B2(data_w[3]), 
        .ZN(n2408) );
  INV_X1 U4036 ( .A(n2409), .ZN(n8796) );
  AOI22_X1 U4037 ( .A1(reg_mem[76]), .A2(n2405), .B1(n8800), .B2(data_w[4]), 
        .ZN(n2409) );
  INV_X1 U4038 ( .A(n2410), .ZN(n8797) );
  AOI22_X1 U4039 ( .A1(reg_mem[77]), .A2(n2405), .B1(n8800), .B2(data_w[5]), 
        .ZN(n2410) );
  INV_X1 U4040 ( .A(n2411), .ZN(n8798) );
  AOI22_X1 U4041 ( .A1(reg_mem[78]), .A2(n2405), .B1(n8800), .B2(data_w[6]), 
        .ZN(n2411) );
  INV_X1 U4042 ( .A(n2412), .ZN(n8799) );
  AOI22_X1 U4043 ( .A1(reg_mem[79]), .A2(n2405), .B1(n8800), .B2(data_w[7]), 
        .ZN(n2412) );
  INV_X1 U4044 ( .A(n2414), .ZN(n7639) );
  AOI22_X1 U4045 ( .A1(reg_mem[80]), .A2(n2415), .B1(n7647), .B2(data_w[0]), 
        .ZN(n2414) );
  INV_X1 U4046 ( .A(n2416), .ZN(n7640) );
  AOI22_X1 U4047 ( .A1(reg_mem[81]), .A2(n2415), .B1(n7647), .B2(data_w[1]), 
        .ZN(n2416) );
  INV_X1 U4048 ( .A(n2417), .ZN(n7641) );
  AOI22_X1 U4049 ( .A1(reg_mem[82]), .A2(n2415), .B1(n7647), .B2(data_w[2]), 
        .ZN(n2417) );
  INV_X1 U4050 ( .A(n2418), .ZN(n7642) );
  AOI22_X1 U4051 ( .A1(reg_mem[83]), .A2(n2415), .B1(n7647), .B2(data_w[3]), 
        .ZN(n2418) );
  INV_X1 U4052 ( .A(n2419), .ZN(n7643) );
  AOI22_X1 U4053 ( .A1(reg_mem[84]), .A2(n2415), .B1(n7647), .B2(data_w[4]), 
        .ZN(n2419) );
  INV_X1 U4054 ( .A(n2420), .ZN(n7644) );
  AOI22_X1 U4055 ( .A1(reg_mem[85]), .A2(n2415), .B1(n7647), .B2(data_w[5]), 
        .ZN(n2420) );
  INV_X1 U4056 ( .A(n2421), .ZN(n7645) );
  AOI22_X1 U4057 ( .A1(reg_mem[86]), .A2(n2415), .B1(n7647), .B2(data_w[6]), 
        .ZN(n2421) );
  INV_X1 U4058 ( .A(n2422), .ZN(n7646) );
  AOI22_X1 U4059 ( .A1(reg_mem[87]), .A2(n2415), .B1(n7647), .B2(data_w[7]), 
        .ZN(n2422) );
  INV_X1 U4060 ( .A(n2424), .ZN(n8216) );
  AOI22_X1 U4061 ( .A1(reg_mem[88]), .A2(n2425), .B1(n8224), .B2(data_w[0]), 
        .ZN(n2424) );
  INV_X1 U4062 ( .A(n2426), .ZN(n8217) );
  AOI22_X1 U4063 ( .A1(reg_mem[89]), .A2(n2425), .B1(n8224), .B2(data_w[1]), 
        .ZN(n2426) );
  INV_X1 U4064 ( .A(n2427), .ZN(n8218) );
  AOI22_X1 U4065 ( .A1(reg_mem[90]), .A2(n2425), .B1(n8224), .B2(data_w[2]), 
        .ZN(n2427) );
  INV_X1 U4066 ( .A(n2428), .ZN(n8219) );
  AOI22_X1 U4067 ( .A1(reg_mem[91]), .A2(n2425), .B1(n8224), .B2(data_w[3]), 
        .ZN(n2428) );
  INV_X1 U4068 ( .A(n2429), .ZN(n8220) );
  AOI22_X1 U4069 ( .A1(reg_mem[92]), .A2(n2425), .B1(n8224), .B2(data_w[4]), 
        .ZN(n2429) );
  INV_X1 U4070 ( .A(n2430), .ZN(n8221) );
  AOI22_X1 U4071 ( .A1(reg_mem[93]), .A2(n2425), .B1(n8224), .B2(data_w[5]), 
        .ZN(n2430) );
  INV_X1 U4072 ( .A(n2431), .ZN(n8222) );
  AOI22_X1 U4073 ( .A1(reg_mem[94]), .A2(n2425), .B1(n8224), .B2(data_w[6]), 
        .ZN(n2431) );
  INV_X1 U4074 ( .A(n2432), .ZN(n8223) );
  AOI22_X1 U4075 ( .A1(reg_mem[95]), .A2(n2425), .B1(n8224), .B2(data_w[7]), 
        .ZN(n2432) );
  INV_X1 U4076 ( .A(n2434), .ZN(n6919) );
  AOI22_X1 U4077 ( .A1(reg_mem[96]), .A2(n2435), .B1(n6927), .B2(data_w[0]), 
        .ZN(n2434) );
  INV_X1 U4078 ( .A(n2436), .ZN(n6920) );
  AOI22_X1 U4079 ( .A1(reg_mem[97]), .A2(n2435), .B1(n6927), .B2(data_w[1]), 
        .ZN(n2436) );
  INV_X1 U4080 ( .A(n2437), .ZN(n6921) );
  AOI22_X1 U4081 ( .A1(reg_mem[98]), .A2(n2435), .B1(n6927), .B2(data_w[2]), 
        .ZN(n2437) );
  INV_X1 U4082 ( .A(n2438), .ZN(n6922) );
  AOI22_X1 U4083 ( .A1(reg_mem[99]), .A2(n2435), .B1(n6927), .B2(data_w[3]), 
        .ZN(n2438) );
  INV_X1 U4084 ( .A(n2439), .ZN(n6923) );
  AOI22_X1 U4085 ( .A1(reg_mem[100]), .A2(n2435), .B1(n6927), .B2(data_w[4]), 
        .ZN(n2439) );
  INV_X1 U4086 ( .A(n2440), .ZN(n6924) );
  AOI22_X1 U4087 ( .A1(reg_mem[101]), .A2(n2435), .B1(n6927), .B2(data_w[5]), 
        .ZN(n2440) );
  INV_X1 U4088 ( .A(n2441), .ZN(n6925) );
  AOI22_X1 U4089 ( .A1(reg_mem[102]), .A2(n2435), .B1(n6927), .B2(data_w[6]), 
        .ZN(n2441) );
  INV_X1 U4090 ( .A(n2442), .ZN(n6926) );
  AOI22_X1 U4091 ( .A1(reg_mem[103]), .A2(n2435), .B1(n6927), .B2(data_w[7]), 
        .ZN(n2442) );
  INV_X1 U4092 ( .A(n2444), .ZN(n8648) );
  AOI22_X1 U4093 ( .A1(reg_mem[104]), .A2(n2445), .B1(n8656), .B2(data_w[0]), 
        .ZN(n2444) );
  INV_X1 U4094 ( .A(n2446), .ZN(n8649) );
  AOI22_X1 U4095 ( .A1(reg_mem[105]), .A2(n2445), .B1(n8656), .B2(data_w[1]), 
        .ZN(n2446) );
  INV_X1 U4096 ( .A(n2447), .ZN(n8650) );
  AOI22_X1 U4097 ( .A1(reg_mem[106]), .A2(n2445), .B1(n8656), .B2(data_w[2]), 
        .ZN(n2447) );
  INV_X1 U4098 ( .A(n2448), .ZN(n8651) );
  AOI22_X1 U4099 ( .A1(reg_mem[107]), .A2(n2445), .B1(n8656), .B2(data_w[3]), 
        .ZN(n2448) );
  INV_X1 U4100 ( .A(n2449), .ZN(n8652) );
  AOI22_X1 U4101 ( .A1(reg_mem[108]), .A2(n2445), .B1(n8656), .B2(data_w[4]), 
        .ZN(n2449) );
  INV_X1 U4102 ( .A(n2450), .ZN(n8653) );
  AOI22_X1 U4103 ( .A1(reg_mem[109]), .A2(n2445), .B1(n8656), .B2(data_w[5]), 
        .ZN(n2450) );
  INV_X1 U4104 ( .A(n2451), .ZN(n8654) );
  AOI22_X1 U4105 ( .A1(reg_mem[110]), .A2(n2445), .B1(n8656), .B2(data_w[6]), 
        .ZN(n2451) );
  INV_X1 U4106 ( .A(n2452), .ZN(n8655) );
  AOI22_X1 U4107 ( .A1(reg_mem[111]), .A2(n2445), .B1(n8656), .B2(data_w[7]), 
        .ZN(n2452) );
  INV_X1 U4108 ( .A(n2454), .ZN(n7495) );
  AOI22_X1 U4109 ( .A1(reg_mem[112]), .A2(n2455), .B1(n7503), .B2(data_w[0]), 
        .ZN(n2454) );
  INV_X1 U4110 ( .A(n2456), .ZN(n7496) );
  AOI22_X1 U4111 ( .A1(reg_mem[113]), .A2(n2455), .B1(n7503), .B2(data_w[1]), 
        .ZN(n2456) );
  INV_X1 U4112 ( .A(n2457), .ZN(n7497) );
  AOI22_X1 U4113 ( .A1(reg_mem[114]), .A2(n2455), .B1(n7503), .B2(data_w[2]), 
        .ZN(n2457) );
  INV_X1 U4114 ( .A(n2458), .ZN(n7498) );
  AOI22_X1 U4115 ( .A1(reg_mem[115]), .A2(n2455), .B1(n7503), .B2(data_w[3]), 
        .ZN(n2458) );
  INV_X1 U4116 ( .A(n2459), .ZN(n7499) );
  AOI22_X1 U4117 ( .A1(reg_mem[116]), .A2(n2455), .B1(n7503), .B2(data_w[4]), 
        .ZN(n2459) );
  INV_X1 U4118 ( .A(n2460), .ZN(n7500) );
  AOI22_X1 U4119 ( .A1(reg_mem[117]), .A2(n2455), .B1(n7503), .B2(data_w[5]), 
        .ZN(n2460) );
  INV_X1 U4120 ( .A(n2461), .ZN(n7501) );
  AOI22_X1 U4121 ( .A1(reg_mem[118]), .A2(n2455), .B1(n7503), .B2(data_w[6]), 
        .ZN(n2461) );
  INV_X1 U4122 ( .A(n2462), .ZN(n7502) );
  AOI22_X1 U4123 ( .A1(reg_mem[119]), .A2(n2455), .B1(n7503), .B2(data_w[7]), 
        .ZN(n2462) );
  INV_X1 U4124 ( .A(n2464), .ZN(n8072) );
  AOI22_X1 U4125 ( .A1(reg_mem[120]), .A2(n2465), .B1(n8080), .B2(data_w[0]), 
        .ZN(n2464) );
  INV_X1 U4126 ( .A(n2466), .ZN(n8073) );
  AOI22_X1 U4127 ( .A1(reg_mem[121]), .A2(n2465), .B1(n8080), .B2(data_w[1]), 
        .ZN(n2466) );
  INV_X1 U4128 ( .A(n2467), .ZN(n8074) );
  AOI22_X1 U4129 ( .A1(reg_mem[122]), .A2(n2465), .B1(n8080), .B2(data_w[2]), 
        .ZN(n2467) );
  INV_X1 U4130 ( .A(n2468), .ZN(n8075) );
  AOI22_X1 U4131 ( .A1(reg_mem[123]), .A2(n2465), .B1(n8080), .B2(data_w[3]), 
        .ZN(n2468) );
  INV_X1 U4132 ( .A(n2469), .ZN(n8076) );
  AOI22_X1 U4133 ( .A1(reg_mem[124]), .A2(n2465), .B1(n8080), .B2(data_w[4]), 
        .ZN(n2469) );
  INV_X1 U4134 ( .A(n2470), .ZN(n8077) );
  AOI22_X1 U4135 ( .A1(reg_mem[125]), .A2(n2465), .B1(n8080), .B2(data_w[5]), 
        .ZN(n2470) );
  INV_X1 U4136 ( .A(n2471), .ZN(n8078) );
  AOI22_X1 U4137 ( .A1(reg_mem[126]), .A2(n2465), .B1(n8080), .B2(data_w[6]), 
        .ZN(n2471) );
  INV_X1 U4138 ( .A(n2472), .ZN(n8079) );
  AOI22_X1 U4139 ( .A1(reg_mem[127]), .A2(n2465), .B1(n8080), .B2(data_w[7]), 
        .ZN(n2472) );
  INV_X1 U4140 ( .A(n2476), .ZN(n7342) );
  AOI22_X1 U4141 ( .A1(reg_mem[128]), .A2(n2477), .B1(n7350), .B2(data_w[0]), 
        .ZN(n2476) );
  INV_X1 U4142 ( .A(n2478), .ZN(n7343) );
  AOI22_X1 U4143 ( .A1(reg_mem[129]), .A2(n2477), .B1(n7350), .B2(data_w[1]), 
        .ZN(n2478) );
  INV_X1 U4144 ( .A(n2479), .ZN(n7344) );
  AOI22_X1 U4145 ( .A1(reg_mem[130]), .A2(n2477), .B1(n7350), .B2(data_w[2]), 
        .ZN(n2479) );
  INV_X1 U4146 ( .A(n2480), .ZN(n7345) );
  AOI22_X1 U4147 ( .A1(reg_mem[131]), .A2(n2477), .B1(n7350), .B2(data_w[3]), 
        .ZN(n2480) );
  INV_X1 U4148 ( .A(n2481), .ZN(n7346) );
  AOI22_X1 U4149 ( .A1(reg_mem[132]), .A2(n2477), .B1(n7350), .B2(data_w[4]), 
        .ZN(n2481) );
  INV_X1 U4150 ( .A(n2482), .ZN(n7347) );
  AOI22_X1 U4151 ( .A1(reg_mem[133]), .A2(n2477), .B1(n7350), .B2(data_w[5]), 
        .ZN(n2482) );
  INV_X1 U4152 ( .A(n2483), .ZN(n7348) );
  AOI22_X1 U4153 ( .A1(reg_mem[134]), .A2(n2477), .B1(n7350), .B2(data_w[6]), 
        .ZN(n2483) );
  INV_X1 U4154 ( .A(n2484), .ZN(n7349) );
  AOI22_X1 U4155 ( .A1(reg_mem[135]), .A2(n2477), .B1(n7350), .B2(data_w[7]), 
        .ZN(n2484) );
  INV_X1 U4156 ( .A(n2486), .ZN(n9071) );
  AOI22_X1 U4157 ( .A1(reg_mem[136]), .A2(n2487), .B1(n9079), .B2(data_w[0]), 
        .ZN(n2486) );
  INV_X1 U4158 ( .A(n2488), .ZN(n9072) );
  AOI22_X1 U4159 ( .A1(reg_mem[137]), .A2(n2487), .B1(n9079), .B2(data_w[1]), 
        .ZN(n2488) );
  INV_X1 U4160 ( .A(n2489), .ZN(n9073) );
  AOI22_X1 U4161 ( .A1(reg_mem[138]), .A2(n2487), .B1(n9079), .B2(data_w[2]), 
        .ZN(n2489) );
  INV_X1 U4162 ( .A(n2490), .ZN(n9074) );
  AOI22_X1 U4163 ( .A1(reg_mem[139]), .A2(n2487), .B1(n9079), .B2(data_w[3]), 
        .ZN(n2490) );
  INV_X1 U4164 ( .A(n2491), .ZN(n9075) );
  AOI22_X1 U4165 ( .A1(reg_mem[140]), .A2(n2487), .B1(n9079), .B2(data_w[4]), 
        .ZN(n2491) );
  INV_X1 U4166 ( .A(n2492), .ZN(n9076) );
  AOI22_X1 U4167 ( .A1(reg_mem[141]), .A2(n2487), .B1(n9079), .B2(data_w[5]), 
        .ZN(n2492) );
  INV_X1 U4168 ( .A(n2493), .ZN(n9077) );
  AOI22_X1 U4169 ( .A1(reg_mem[142]), .A2(n2487), .B1(n9079), .B2(data_w[6]), 
        .ZN(n2493) );
  INV_X1 U4170 ( .A(n2494), .ZN(n9078) );
  AOI22_X1 U4171 ( .A1(reg_mem[143]), .A2(n2487), .B1(n9079), .B2(data_w[7]), 
        .ZN(n2494) );
  INV_X1 U4172 ( .A(n2495), .ZN(n7918) );
  AOI22_X1 U4173 ( .A1(reg_mem[144]), .A2(n2496), .B1(n7926), .B2(data_w[0]), 
        .ZN(n2495) );
  INV_X1 U4174 ( .A(n2497), .ZN(n7919) );
  AOI22_X1 U4175 ( .A1(reg_mem[145]), .A2(n2496), .B1(n7926), .B2(data_w[1]), 
        .ZN(n2497) );
  INV_X1 U4176 ( .A(n2498), .ZN(n7920) );
  AOI22_X1 U4177 ( .A1(reg_mem[146]), .A2(n2496), .B1(n7926), .B2(data_w[2]), 
        .ZN(n2498) );
  INV_X1 U4178 ( .A(n2499), .ZN(n7921) );
  AOI22_X1 U4179 ( .A1(reg_mem[147]), .A2(n2496), .B1(n7926), .B2(data_w[3]), 
        .ZN(n2499) );
  INV_X1 U4180 ( .A(n2500), .ZN(n7922) );
  AOI22_X1 U4181 ( .A1(reg_mem[148]), .A2(n2496), .B1(n7926), .B2(data_w[4]), 
        .ZN(n2500) );
  INV_X1 U4182 ( .A(n2501), .ZN(n7923) );
  AOI22_X1 U4183 ( .A1(reg_mem[149]), .A2(n2496), .B1(n7926), .B2(data_w[5]), 
        .ZN(n2501) );
  INV_X1 U4184 ( .A(n2502), .ZN(n7924) );
  AOI22_X1 U4185 ( .A1(reg_mem[150]), .A2(n2496), .B1(n7926), .B2(data_w[6]), 
        .ZN(n2502) );
  INV_X1 U4186 ( .A(n2503), .ZN(n7925) );
  AOI22_X1 U4187 ( .A1(reg_mem[151]), .A2(n2496), .B1(n7926), .B2(data_w[7]), 
        .ZN(n2503) );
  INV_X1 U4188 ( .A(n2504), .ZN(n8495) );
  AOI22_X1 U4189 ( .A1(reg_mem[152]), .A2(n2505), .B1(n8503), .B2(data_w[0]), 
        .ZN(n2504) );
  INV_X1 U4190 ( .A(n2506), .ZN(n8496) );
  AOI22_X1 U4191 ( .A1(reg_mem[153]), .A2(n2505), .B1(n8503), .B2(data_w[1]), 
        .ZN(n2506) );
  INV_X1 U4192 ( .A(n2507), .ZN(n8497) );
  AOI22_X1 U4193 ( .A1(reg_mem[154]), .A2(n2505), .B1(n8503), .B2(data_w[2]), 
        .ZN(n2507) );
  INV_X1 U4194 ( .A(n2508), .ZN(n8498) );
  AOI22_X1 U4195 ( .A1(reg_mem[155]), .A2(n2505), .B1(n8503), .B2(data_w[3]), 
        .ZN(n2508) );
  INV_X1 U4196 ( .A(n2509), .ZN(n8499) );
  AOI22_X1 U4197 ( .A1(reg_mem[156]), .A2(n2505), .B1(n8503), .B2(data_w[4]), 
        .ZN(n2509) );
  INV_X1 U4198 ( .A(n2510), .ZN(n8500) );
  AOI22_X1 U4199 ( .A1(reg_mem[157]), .A2(n2505), .B1(n8503), .B2(data_w[5]), 
        .ZN(n2510) );
  INV_X1 U4200 ( .A(n2511), .ZN(n8501) );
  AOI22_X1 U4201 ( .A1(reg_mem[158]), .A2(n2505), .B1(n8503), .B2(data_w[6]), 
        .ZN(n2511) );
  INV_X1 U4202 ( .A(n2512), .ZN(n8502) );
  AOI22_X1 U4203 ( .A1(reg_mem[159]), .A2(n2505), .B1(n8503), .B2(data_w[7]), 
        .ZN(n2512) );
  INV_X1 U4204 ( .A(n2513), .ZN(n7198) );
  AOI22_X1 U4205 ( .A1(reg_mem[160]), .A2(n2514), .B1(n7206), .B2(data_w[0]), 
        .ZN(n2513) );
  INV_X1 U4206 ( .A(n2515), .ZN(n7199) );
  AOI22_X1 U4207 ( .A1(reg_mem[161]), .A2(n2514), .B1(n7206), .B2(data_w[1]), 
        .ZN(n2515) );
  INV_X1 U4208 ( .A(n2516), .ZN(n7200) );
  AOI22_X1 U4209 ( .A1(reg_mem[162]), .A2(n2514), .B1(n7206), .B2(data_w[2]), 
        .ZN(n2516) );
  INV_X1 U4210 ( .A(n2517), .ZN(n7201) );
  AOI22_X1 U4211 ( .A1(reg_mem[163]), .A2(n2514), .B1(n7206), .B2(data_w[3]), 
        .ZN(n2517) );
  INV_X1 U4212 ( .A(n2518), .ZN(n7202) );
  AOI22_X1 U4213 ( .A1(reg_mem[164]), .A2(n2514), .B1(n7206), .B2(data_w[4]), 
        .ZN(n2518) );
  INV_X1 U4214 ( .A(n2519), .ZN(n7203) );
  AOI22_X1 U4215 ( .A1(reg_mem[165]), .A2(n2514), .B1(n7206), .B2(data_w[5]), 
        .ZN(n2519) );
  INV_X1 U4216 ( .A(n2520), .ZN(n7204) );
  AOI22_X1 U4217 ( .A1(reg_mem[166]), .A2(n2514), .B1(n7206), .B2(data_w[6]), 
        .ZN(n2520) );
  INV_X1 U4218 ( .A(n2521), .ZN(n7205) );
  AOI22_X1 U4219 ( .A1(reg_mem[167]), .A2(n2514), .B1(n7206), .B2(data_w[7]), 
        .ZN(n2521) );
  INV_X1 U4220 ( .A(n2522), .ZN(n8927) );
  AOI22_X1 U4221 ( .A1(reg_mem[168]), .A2(n2523), .B1(n8935), .B2(data_w[0]), 
        .ZN(n2522) );
  INV_X1 U4222 ( .A(n2524), .ZN(n8928) );
  AOI22_X1 U4223 ( .A1(reg_mem[169]), .A2(n2523), .B1(n8935), .B2(data_w[1]), 
        .ZN(n2524) );
  INV_X1 U4224 ( .A(n2525), .ZN(n8929) );
  AOI22_X1 U4225 ( .A1(reg_mem[170]), .A2(n2523), .B1(n8935), .B2(data_w[2]), 
        .ZN(n2525) );
  INV_X1 U4226 ( .A(n2526), .ZN(n8930) );
  AOI22_X1 U4227 ( .A1(reg_mem[171]), .A2(n2523), .B1(n8935), .B2(data_w[3]), 
        .ZN(n2526) );
  INV_X1 U4228 ( .A(n2527), .ZN(n8931) );
  AOI22_X1 U4229 ( .A1(reg_mem[172]), .A2(n2523), .B1(n8935), .B2(data_w[4]), 
        .ZN(n2527) );
  INV_X1 U4230 ( .A(n2528), .ZN(n8932) );
  AOI22_X1 U4231 ( .A1(reg_mem[173]), .A2(n2523), .B1(n8935), .B2(data_w[5]), 
        .ZN(n2528) );
  INV_X1 U4232 ( .A(n2529), .ZN(n8933) );
  AOI22_X1 U4233 ( .A1(reg_mem[174]), .A2(n2523), .B1(n8935), .B2(data_w[6]), 
        .ZN(n2529) );
  INV_X1 U4234 ( .A(n2530), .ZN(n8934) );
  AOI22_X1 U4235 ( .A1(reg_mem[175]), .A2(n2523), .B1(n8935), .B2(data_w[7]), 
        .ZN(n2530) );
  INV_X1 U4236 ( .A(n2531), .ZN(n7774) );
  AOI22_X1 U4237 ( .A1(reg_mem[176]), .A2(n2532), .B1(n7782), .B2(data_w[0]), 
        .ZN(n2531) );
  INV_X1 U4238 ( .A(n2533), .ZN(n7775) );
  AOI22_X1 U4239 ( .A1(reg_mem[177]), .A2(n2532), .B1(n7782), .B2(data_w[1]), 
        .ZN(n2533) );
  INV_X1 U4240 ( .A(n2534), .ZN(n7776) );
  AOI22_X1 U4241 ( .A1(reg_mem[178]), .A2(n2532), .B1(n7782), .B2(data_w[2]), 
        .ZN(n2534) );
  INV_X1 U4242 ( .A(n2535), .ZN(n7777) );
  AOI22_X1 U4243 ( .A1(reg_mem[179]), .A2(n2532), .B1(n7782), .B2(data_w[3]), 
        .ZN(n2535) );
  INV_X1 U4244 ( .A(n2536), .ZN(n7778) );
  AOI22_X1 U4245 ( .A1(reg_mem[180]), .A2(n2532), .B1(n7782), .B2(data_w[4]), 
        .ZN(n2536) );
  INV_X1 U4246 ( .A(n2537), .ZN(n7779) );
  AOI22_X1 U4247 ( .A1(reg_mem[181]), .A2(n2532), .B1(n7782), .B2(data_w[5]), 
        .ZN(n2537) );
  INV_X1 U4248 ( .A(n2538), .ZN(n7780) );
  AOI22_X1 U4249 ( .A1(reg_mem[182]), .A2(n2532), .B1(n7782), .B2(data_w[6]), 
        .ZN(n2538) );
  INV_X1 U4250 ( .A(n2539), .ZN(n7781) );
  AOI22_X1 U4251 ( .A1(reg_mem[183]), .A2(n2532), .B1(n7782), .B2(data_w[7]), 
        .ZN(n2539) );
  INV_X1 U4252 ( .A(n2540), .ZN(n8351) );
  AOI22_X1 U4253 ( .A1(reg_mem[184]), .A2(n2541), .B1(n8359), .B2(data_w[0]), 
        .ZN(n2540) );
  INV_X1 U4254 ( .A(n2542), .ZN(n8352) );
  AOI22_X1 U4255 ( .A1(reg_mem[185]), .A2(n2541), .B1(n8359), .B2(data_w[1]), 
        .ZN(n2542) );
  INV_X1 U4256 ( .A(n2543), .ZN(n8353) );
  AOI22_X1 U4257 ( .A1(reg_mem[186]), .A2(n2541), .B1(n8359), .B2(data_w[2]), 
        .ZN(n2543) );
  INV_X1 U4258 ( .A(n2544), .ZN(n8354) );
  AOI22_X1 U4259 ( .A1(reg_mem[187]), .A2(n2541), .B1(n8359), .B2(data_w[3]), 
        .ZN(n2544) );
  INV_X1 U4260 ( .A(n2545), .ZN(n8355) );
  AOI22_X1 U4261 ( .A1(reg_mem[188]), .A2(n2541), .B1(n8359), .B2(data_w[4]), 
        .ZN(n2545) );
  INV_X1 U4262 ( .A(n2546), .ZN(n8356) );
  AOI22_X1 U4263 ( .A1(reg_mem[189]), .A2(n2541), .B1(n8359), .B2(data_w[5]), 
        .ZN(n2546) );
  INV_X1 U4264 ( .A(n2547), .ZN(n8357) );
  AOI22_X1 U4265 ( .A1(reg_mem[190]), .A2(n2541), .B1(n8359), .B2(data_w[6]), 
        .ZN(n2547) );
  INV_X1 U4266 ( .A(n2548), .ZN(n8358) );
  AOI22_X1 U4267 ( .A1(reg_mem[191]), .A2(n2541), .B1(n8359), .B2(data_w[7]), 
        .ZN(n2548) );
  INV_X1 U4268 ( .A(n2549), .ZN(n7054) );
  AOI22_X1 U4269 ( .A1(reg_mem[192]), .A2(n2550), .B1(n7062), .B2(data_w[0]), 
        .ZN(n2549) );
  INV_X1 U4270 ( .A(n2551), .ZN(n7055) );
  AOI22_X1 U4271 ( .A1(reg_mem[193]), .A2(n2550), .B1(n7062), .B2(data_w[1]), 
        .ZN(n2551) );
  INV_X1 U4272 ( .A(n2552), .ZN(n7056) );
  AOI22_X1 U4273 ( .A1(reg_mem[194]), .A2(n2550), .B1(n7062), .B2(data_w[2]), 
        .ZN(n2552) );
  INV_X1 U4274 ( .A(n2553), .ZN(n7057) );
  AOI22_X1 U4275 ( .A1(reg_mem[195]), .A2(n2550), .B1(n7062), .B2(data_w[3]), 
        .ZN(n2553) );
  INV_X1 U4276 ( .A(n2554), .ZN(n7058) );
  AOI22_X1 U4277 ( .A1(reg_mem[196]), .A2(n2550), .B1(n7062), .B2(data_w[4]), 
        .ZN(n2554) );
  INV_X1 U4278 ( .A(n2555), .ZN(n7059) );
  AOI22_X1 U4279 ( .A1(reg_mem[197]), .A2(n2550), .B1(n7062), .B2(data_w[5]), 
        .ZN(n2555) );
  INV_X1 U4280 ( .A(n2556), .ZN(n7060) );
  AOI22_X1 U4281 ( .A1(reg_mem[198]), .A2(n2550), .B1(n7062), .B2(data_w[6]), 
        .ZN(n2556) );
  INV_X1 U4282 ( .A(n2557), .ZN(n7061) );
  AOI22_X1 U4283 ( .A1(reg_mem[199]), .A2(n2550), .B1(n7062), .B2(data_w[7]), 
        .ZN(n2557) );
  INV_X1 U4284 ( .A(n2558), .ZN(n8783) );
  AOI22_X1 U4285 ( .A1(reg_mem[200]), .A2(n2559), .B1(n8791), .B2(data_w[0]), 
        .ZN(n2558) );
  INV_X1 U4286 ( .A(n2560), .ZN(n8784) );
  AOI22_X1 U4287 ( .A1(reg_mem[201]), .A2(n2559), .B1(n8791), .B2(data_w[1]), 
        .ZN(n2560) );
  INV_X1 U4288 ( .A(n2561), .ZN(n8785) );
  AOI22_X1 U4289 ( .A1(reg_mem[202]), .A2(n2559), .B1(n8791), .B2(data_w[2]), 
        .ZN(n2561) );
  INV_X1 U4290 ( .A(n2562), .ZN(n8786) );
  AOI22_X1 U4291 ( .A1(reg_mem[203]), .A2(n2559), .B1(n8791), .B2(data_w[3]), 
        .ZN(n2562) );
  INV_X1 U4292 ( .A(n2563), .ZN(n8787) );
  AOI22_X1 U4293 ( .A1(reg_mem[204]), .A2(n2559), .B1(n8791), .B2(data_w[4]), 
        .ZN(n2563) );
  INV_X1 U4294 ( .A(n2564), .ZN(n8788) );
  AOI22_X1 U4295 ( .A1(reg_mem[205]), .A2(n2559), .B1(n8791), .B2(data_w[5]), 
        .ZN(n2564) );
  INV_X1 U4296 ( .A(n2565), .ZN(n8789) );
  AOI22_X1 U4297 ( .A1(reg_mem[206]), .A2(n2559), .B1(n8791), .B2(data_w[6]), 
        .ZN(n2565) );
  INV_X1 U4298 ( .A(n2566), .ZN(n8790) );
  AOI22_X1 U4299 ( .A1(reg_mem[207]), .A2(n2559), .B1(n8791), .B2(data_w[7]), 
        .ZN(n2566) );
  INV_X1 U4300 ( .A(n2567), .ZN(n7630) );
  AOI22_X1 U4301 ( .A1(reg_mem[208]), .A2(n2568), .B1(n7638), .B2(data_w[0]), 
        .ZN(n2567) );
  INV_X1 U4302 ( .A(n2569), .ZN(n7631) );
  AOI22_X1 U4303 ( .A1(reg_mem[209]), .A2(n2568), .B1(n7638), .B2(data_w[1]), 
        .ZN(n2569) );
  INV_X1 U4304 ( .A(n2570), .ZN(n7632) );
  AOI22_X1 U4305 ( .A1(reg_mem[210]), .A2(n2568), .B1(n7638), .B2(data_w[2]), 
        .ZN(n2570) );
  INV_X1 U4306 ( .A(n2571), .ZN(n7633) );
  AOI22_X1 U4307 ( .A1(reg_mem[211]), .A2(n2568), .B1(n7638), .B2(data_w[3]), 
        .ZN(n2571) );
  INV_X1 U4308 ( .A(n2572), .ZN(n7634) );
  AOI22_X1 U4309 ( .A1(reg_mem[212]), .A2(n2568), .B1(n7638), .B2(data_w[4]), 
        .ZN(n2572) );
  INV_X1 U4310 ( .A(n2573), .ZN(n7635) );
  AOI22_X1 U4311 ( .A1(reg_mem[213]), .A2(n2568), .B1(n7638), .B2(data_w[5]), 
        .ZN(n2573) );
  INV_X1 U4312 ( .A(n2574), .ZN(n7636) );
  AOI22_X1 U4313 ( .A1(reg_mem[214]), .A2(n2568), .B1(n7638), .B2(data_w[6]), 
        .ZN(n2574) );
  INV_X1 U4314 ( .A(n2575), .ZN(n7637) );
  AOI22_X1 U4315 ( .A1(reg_mem[215]), .A2(n2568), .B1(n7638), .B2(data_w[7]), 
        .ZN(n2575) );
  INV_X1 U4316 ( .A(n2576), .ZN(n8207) );
  AOI22_X1 U4317 ( .A1(reg_mem[216]), .A2(n2577), .B1(n8215), .B2(data_w[0]), 
        .ZN(n2576) );
  INV_X1 U4318 ( .A(n2578), .ZN(n8208) );
  AOI22_X1 U4319 ( .A1(reg_mem[217]), .A2(n2577), .B1(n8215), .B2(data_w[1]), 
        .ZN(n2578) );
  INV_X1 U4320 ( .A(n2579), .ZN(n8209) );
  AOI22_X1 U4321 ( .A1(reg_mem[218]), .A2(n2577), .B1(n8215), .B2(data_w[2]), 
        .ZN(n2579) );
  INV_X1 U4322 ( .A(n2580), .ZN(n8210) );
  AOI22_X1 U4323 ( .A1(reg_mem[219]), .A2(n2577), .B1(n8215), .B2(data_w[3]), 
        .ZN(n2580) );
  INV_X1 U4324 ( .A(n2581), .ZN(n8211) );
  AOI22_X1 U4325 ( .A1(reg_mem[220]), .A2(n2577), .B1(n8215), .B2(data_w[4]), 
        .ZN(n2581) );
  INV_X1 U4326 ( .A(n2582), .ZN(n8212) );
  AOI22_X1 U4327 ( .A1(reg_mem[221]), .A2(n2577), .B1(n8215), .B2(data_w[5]), 
        .ZN(n2582) );
  INV_X1 U4328 ( .A(n2583), .ZN(n8213) );
  AOI22_X1 U4329 ( .A1(reg_mem[222]), .A2(n2577), .B1(n8215), .B2(data_w[6]), 
        .ZN(n2583) );
  INV_X1 U4330 ( .A(n2584), .ZN(n8214) );
  AOI22_X1 U4331 ( .A1(reg_mem[223]), .A2(n2577), .B1(n8215), .B2(data_w[7]), 
        .ZN(n2584) );
  INV_X1 U4332 ( .A(n2585), .ZN(n6910) );
  AOI22_X1 U4333 ( .A1(reg_mem[224]), .A2(n2586), .B1(n6918), .B2(data_w[0]), 
        .ZN(n2585) );
  INV_X1 U4334 ( .A(n2587), .ZN(n6911) );
  AOI22_X1 U4335 ( .A1(reg_mem[225]), .A2(n2586), .B1(n6918), .B2(data_w[1]), 
        .ZN(n2587) );
  INV_X1 U4336 ( .A(n2588), .ZN(n6912) );
  AOI22_X1 U4337 ( .A1(reg_mem[226]), .A2(n2586), .B1(n6918), .B2(data_w[2]), 
        .ZN(n2588) );
  INV_X1 U4338 ( .A(n2589), .ZN(n6913) );
  AOI22_X1 U4339 ( .A1(reg_mem[227]), .A2(n2586), .B1(n6918), .B2(data_w[3]), 
        .ZN(n2589) );
  INV_X1 U4340 ( .A(n2590), .ZN(n6914) );
  AOI22_X1 U4341 ( .A1(reg_mem[228]), .A2(n2586), .B1(n6918), .B2(data_w[4]), 
        .ZN(n2590) );
  INV_X1 U4342 ( .A(n2591), .ZN(n6915) );
  AOI22_X1 U4343 ( .A1(reg_mem[229]), .A2(n2586), .B1(n6918), .B2(data_w[5]), 
        .ZN(n2591) );
  INV_X1 U4344 ( .A(n2592), .ZN(n6916) );
  AOI22_X1 U4345 ( .A1(reg_mem[230]), .A2(n2586), .B1(n6918), .B2(data_w[6]), 
        .ZN(n2592) );
  INV_X1 U4346 ( .A(n2593), .ZN(n6917) );
  AOI22_X1 U4347 ( .A1(reg_mem[231]), .A2(n2586), .B1(n6918), .B2(data_w[7]), 
        .ZN(n2593) );
  INV_X1 U4348 ( .A(n2594), .ZN(n8639) );
  AOI22_X1 U4349 ( .A1(reg_mem[232]), .A2(n2595), .B1(n8647), .B2(data_w[0]), 
        .ZN(n2594) );
  INV_X1 U4350 ( .A(n2596), .ZN(n8640) );
  AOI22_X1 U4351 ( .A1(reg_mem[233]), .A2(n2595), .B1(n8647), .B2(data_w[1]), 
        .ZN(n2596) );
  INV_X1 U4352 ( .A(n2597), .ZN(n8641) );
  AOI22_X1 U4353 ( .A1(reg_mem[234]), .A2(n2595), .B1(n8647), .B2(data_w[2]), 
        .ZN(n2597) );
  INV_X1 U4354 ( .A(n2598), .ZN(n8642) );
  AOI22_X1 U4355 ( .A1(reg_mem[235]), .A2(n2595), .B1(n8647), .B2(data_w[3]), 
        .ZN(n2598) );
  INV_X1 U4356 ( .A(n2599), .ZN(n8643) );
  AOI22_X1 U4357 ( .A1(reg_mem[236]), .A2(n2595), .B1(n8647), .B2(data_w[4]), 
        .ZN(n2599) );
  INV_X1 U4358 ( .A(n2600), .ZN(n8644) );
  AOI22_X1 U4359 ( .A1(reg_mem[237]), .A2(n2595), .B1(n8647), .B2(data_w[5]), 
        .ZN(n2600) );
  INV_X1 U4360 ( .A(n2601), .ZN(n8645) );
  AOI22_X1 U4361 ( .A1(reg_mem[238]), .A2(n2595), .B1(n8647), .B2(data_w[6]), 
        .ZN(n2601) );
  INV_X1 U4362 ( .A(n2602), .ZN(n8646) );
  AOI22_X1 U4363 ( .A1(reg_mem[239]), .A2(n2595), .B1(n8647), .B2(data_w[7]), 
        .ZN(n2602) );
  INV_X1 U4364 ( .A(n2603), .ZN(n7486) );
  AOI22_X1 U4365 ( .A1(reg_mem[240]), .A2(n2604), .B1(n7494), .B2(data_w[0]), 
        .ZN(n2603) );
  INV_X1 U4366 ( .A(n2605), .ZN(n7487) );
  AOI22_X1 U4367 ( .A1(reg_mem[241]), .A2(n2604), .B1(n7494), .B2(data_w[1]), 
        .ZN(n2605) );
  INV_X1 U4368 ( .A(n2606), .ZN(n7488) );
  AOI22_X1 U4369 ( .A1(reg_mem[242]), .A2(n2604), .B1(n7494), .B2(data_w[2]), 
        .ZN(n2606) );
  INV_X1 U4370 ( .A(n2607), .ZN(n7489) );
  AOI22_X1 U4371 ( .A1(reg_mem[243]), .A2(n2604), .B1(n7494), .B2(data_w[3]), 
        .ZN(n2607) );
  INV_X1 U4372 ( .A(n2608), .ZN(n7490) );
  AOI22_X1 U4373 ( .A1(reg_mem[244]), .A2(n2604), .B1(n7494), .B2(data_w[4]), 
        .ZN(n2608) );
  INV_X1 U4374 ( .A(n2609), .ZN(n7491) );
  AOI22_X1 U4375 ( .A1(reg_mem[245]), .A2(n2604), .B1(n7494), .B2(data_w[5]), 
        .ZN(n2609) );
  INV_X1 U4376 ( .A(n2610), .ZN(n7492) );
  AOI22_X1 U4377 ( .A1(reg_mem[246]), .A2(n2604), .B1(n7494), .B2(data_w[6]), 
        .ZN(n2610) );
  INV_X1 U4378 ( .A(n2611), .ZN(n7493) );
  AOI22_X1 U4379 ( .A1(reg_mem[247]), .A2(n2604), .B1(n7494), .B2(data_w[7]), 
        .ZN(n2611) );
  INV_X1 U4380 ( .A(n2612), .ZN(n8063) );
  AOI22_X1 U4381 ( .A1(reg_mem[248]), .A2(n2613), .B1(n8071), .B2(data_w[0]), 
        .ZN(n2612) );
  INV_X1 U4382 ( .A(n2614), .ZN(n8064) );
  AOI22_X1 U4383 ( .A1(reg_mem[249]), .A2(n2613), .B1(n8071), .B2(data_w[1]), 
        .ZN(n2614) );
  INV_X1 U4384 ( .A(n2615), .ZN(n8065) );
  AOI22_X1 U4385 ( .A1(reg_mem[250]), .A2(n2613), .B1(n8071), .B2(data_w[2]), 
        .ZN(n2615) );
  INV_X1 U4386 ( .A(n2616), .ZN(n8066) );
  AOI22_X1 U4387 ( .A1(reg_mem[251]), .A2(n2613), .B1(n8071), .B2(data_w[3]), 
        .ZN(n2616) );
  INV_X1 U4388 ( .A(n2617), .ZN(n8067) );
  AOI22_X1 U4389 ( .A1(reg_mem[252]), .A2(n2613), .B1(n8071), .B2(data_w[4]), 
        .ZN(n2617) );
  INV_X1 U4390 ( .A(n2618), .ZN(n8068) );
  AOI22_X1 U4391 ( .A1(reg_mem[253]), .A2(n2613), .B1(n8071), .B2(data_w[5]), 
        .ZN(n2618) );
  INV_X1 U4392 ( .A(n2619), .ZN(n8069) );
  AOI22_X1 U4393 ( .A1(reg_mem[254]), .A2(n2613), .B1(n8071), .B2(data_w[6]), 
        .ZN(n2619) );
  INV_X1 U4394 ( .A(n2620), .ZN(n8070) );
  AOI22_X1 U4395 ( .A1(reg_mem[255]), .A2(n2613), .B1(n8071), .B2(data_w[7]), 
        .ZN(n2620) );
  INV_X1 U4396 ( .A(n2622), .ZN(n7333) );
  AOI22_X1 U4397 ( .A1(reg_mem[256]), .A2(n2623), .B1(n7341), .B2(data_w[0]), 
        .ZN(n2622) );
  INV_X1 U4398 ( .A(n2624), .ZN(n7334) );
  AOI22_X1 U4399 ( .A1(reg_mem[257]), .A2(n2623), .B1(n7341), .B2(data_w[1]), 
        .ZN(n2624) );
  INV_X1 U4400 ( .A(n2625), .ZN(n7335) );
  AOI22_X1 U4401 ( .A1(reg_mem[258]), .A2(n2623), .B1(n7341), .B2(data_w[2]), 
        .ZN(n2625) );
  INV_X1 U4402 ( .A(n2626), .ZN(n7336) );
  AOI22_X1 U4403 ( .A1(reg_mem[259]), .A2(n2623), .B1(n7341), .B2(data_w[3]), 
        .ZN(n2626) );
  INV_X1 U4404 ( .A(n2627), .ZN(n7337) );
  AOI22_X1 U4405 ( .A1(reg_mem[260]), .A2(n2623), .B1(n7341), .B2(data_w[4]), 
        .ZN(n2627) );
  INV_X1 U4406 ( .A(n2628), .ZN(n7338) );
  AOI22_X1 U4407 ( .A1(reg_mem[261]), .A2(n2623), .B1(n7341), .B2(data_w[5]), 
        .ZN(n2628) );
  INV_X1 U4408 ( .A(n2629), .ZN(n7339) );
  AOI22_X1 U4409 ( .A1(reg_mem[262]), .A2(n2623), .B1(n7341), .B2(data_w[6]), 
        .ZN(n2629) );
  INV_X1 U4410 ( .A(n2630), .ZN(n7340) );
  AOI22_X1 U4411 ( .A1(reg_mem[263]), .A2(n2623), .B1(n7341), .B2(data_w[7]), 
        .ZN(n2630) );
  INV_X1 U4412 ( .A(n2632), .ZN(n9062) );
  AOI22_X1 U4413 ( .A1(reg_mem[264]), .A2(n2633), .B1(n9070), .B2(data_w[0]), 
        .ZN(n2632) );
  INV_X1 U4414 ( .A(n2634), .ZN(n9063) );
  AOI22_X1 U4415 ( .A1(reg_mem[265]), .A2(n2633), .B1(n9070), .B2(data_w[1]), 
        .ZN(n2634) );
  INV_X1 U4416 ( .A(n2635), .ZN(n9064) );
  AOI22_X1 U4417 ( .A1(reg_mem[266]), .A2(n2633), .B1(n9070), .B2(data_w[2]), 
        .ZN(n2635) );
  INV_X1 U4418 ( .A(n2636), .ZN(n9065) );
  AOI22_X1 U4419 ( .A1(reg_mem[267]), .A2(n2633), .B1(n9070), .B2(data_w[3]), 
        .ZN(n2636) );
  INV_X1 U4420 ( .A(n2637), .ZN(n9066) );
  AOI22_X1 U4421 ( .A1(reg_mem[268]), .A2(n2633), .B1(n9070), .B2(data_w[4]), 
        .ZN(n2637) );
  INV_X1 U4422 ( .A(n2638), .ZN(n9067) );
  AOI22_X1 U4423 ( .A1(reg_mem[269]), .A2(n2633), .B1(n9070), .B2(data_w[5]), 
        .ZN(n2638) );
  INV_X1 U4424 ( .A(n2639), .ZN(n9068) );
  AOI22_X1 U4425 ( .A1(reg_mem[270]), .A2(n2633), .B1(n9070), .B2(data_w[6]), 
        .ZN(n2639) );
  INV_X1 U4426 ( .A(n2640), .ZN(n9069) );
  AOI22_X1 U4427 ( .A1(reg_mem[271]), .A2(n2633), .B1(n9070), .B2(data_w[7]), 
        .ZN(n2640) );
  INV_X1 U4428 ( .A(n2641), .ZN(n7909) );
  AOI22_X1 U4429 ( .A1(reg_mem[272]), .A2(n2642), .B1(n7917), .B2(data_w[0]), 
        .ZN(n2641) );
  INV_X1 U4430 ( .A(n2643), .ZN(n7910) );
  AOI22_X1 U4431 ( .A1(reg_mem[273]), .A2(n2642), .B1(n7917), .B2(data_w[1]), 
        .ZN(n2643) );
  INV_X1 U4432 ( .A(n2644), .ZN(n7911) );
  AOI22_X1 U4433 ( .A1(reg_mem[274]), .A2(n2642), .B1(n7917), .B2(data_w[2]), 
        .ZN(n2644) );
  INV_X1 U4434 ( .A(n2645), .ZN(n7912) );
  AOI22_X1 U4435 ( .A1(reg_mem[275]), .A2(n2642), .B1(n7917), .B2(data_w[3]), 
        .ZN(n2645) );
  INV_X1 U4436 ( .A(n2646), .ZN(n7913) );
  AOI22_X1 U4437 ( .A1(reg_mem[276]), .A2(n2642), .B1(n7917), .B2(data_w[4]), 
        .ZN(n2646) );
  INV_X1 U4438 ( .A(n2647), .ZN(n7914) );
  AOI22_X1 U4439 ( .A1(reg_mem[277]), .A2(n2642), .B1(n7917), .B2(data_w[5]), 
        .ZN(n2647) );
  INV_X1 U4440 ( .A(n2648), .ZN(n7915) );
  AOI22_X1 U4441 ( .A1(reg_mem[278]), .A2(n2642), .B1(n7917), .B2(data_w[6]), 
        .ZN(n2648) );
  INV_X1 U4442 ( .A(n2649), .ZN(n7916) );
  AOI22_X1 U4443 ( .A1(reg_mem[279]), .A2(n2642), .B1(n7917), .B2(data_w[7]), 
        .ZN(n2649) );
  INV_X1 U4444 ( .A(n2650), .ZN(n8486) );
  AOI22_X1 U4445 ( .A1(reg_mem[280]), .A2(n2651), .B1(n8494), .B2(data_w[0]), 
        .ZN(n2650) );
  INV_X1 U4446 ( .A(n2652), .ZN(n8487) );
  AOI22_X1 U4447 ( .A1(reg_mem[281]), .A2(n2651), .B1(n8494), .B2(data_w[1]), 
        .ZN(n2652) );
  INV_X1 U4448 ( .A(n2653), .ZN(n8488) );
  AOI22_X1 U4449 ( .A1(reg_mem[282]), .A2(n2651), .B1(n8494), .B2(data_w[2]), 
        .ZN(n2653) );
  INV_X1 U4450 ( .A(n2654), .ZN(n8489) );
  AOI22_X1 U4451 ( .A1(reg_mem[283]), .A2(n2651), .B1(n8494), .B2(data_w[3]), 
        .ZN(n2654) );
  INV_X1 U4452 ( .A(n2655), .ZN(n8490) );
  AOI22_X1 U4453 ( .A1(reg_mem[284]), .A2(n2651), .B1(n8494), .B2(data_w[4]), 
        .ZN(n2655) );
  INV_X1 U4454 ( .A(n2656), .ZN(n8491) );
  AOI22_X1 U4455 ( .A1(reg_mem[285]), .A2(n2651), .B1(n8494), .B2(data_w[5]), 
        .ZN(n2656) );
  INV_X1 U4456 ( .A(n2657), .ZN(n8492) );
  AOI22_X1 U4457 ( .A1(reg_mem[286]), .A2(n2651), .B1(n8494), .B2(data_w[6]), 
        .ZN(n2657) );
  INV_X1 U4458 ( .A(n2658), .ZN(n8493) );
  AOI22_X1 U4459 ( .A1(reg_mem[287]), .A2(n2651), .B1(n8494), .B2(data_w[7]), 
        .ZN(n2658) );
  INV_X1 U4460 ( .A(n2659), .ZN(n7189) );
  AOI22_X1 U4461 ( .A1(reg_mem[288]), .A2(n2660), .B1(n7197), .B2(data_w[0]), 
        .ZN(n2659) );
  INV_X1 U4462 ( .A(n2661), .ZN(n7190) );
  AOI22_X1 U4463 ( .A1(reg_mem[289]), .A2(n2660), .B1(n7197), .B2(data_w[1]), 
        .ZN(n2661) );
  INV_X1 U4464 ( .A(n2662), .ZN(n7191) );
  AOI22_X1 U4465 ( .A1(reg_mem[290]), .A2(n2660), .B1(n7197), .B2(data_w[2]), 
        .ZN(n2662) );
  INV_X1 U4466 ( .A(n2663), .ZN(n7192) );
  AOI22_X1 U4467 ( .A1(reg_mem[291]), .A2(n2660), .B1(n7197), .B2(data_w[3]), 
        .ZN(n2663) );
  INV_X1 U4468 ( .A(n2664), .ZN(n7193) );
  AOI22_X1 U4469 ( .A1(reg_mem[292]), .A2(n2660), .B1(n7197), .B2(data_w[4]), 
        .ZN(n2664) );
  INV_X1 U4470 ( .A(n2665), .ZN(n7194) );
  AOI22_X1 U4471 ( .A1(reg_mem[293]), .A2(n2660), .B1(n7197), .B2(data_w[5]), 
        .ZN(n2665) );
  INV_X1 U4472 ( .A(n2666), .ZN(n7195) );
  AOI22_X1 U4473 ( .A1(reg_mem[294]), .A2(n2660), .B1(n7197), .B2(data_w[6]), 
        .ZN(n2666) );
  INV_X1 U4474 ( .A(n2667), .ZN(n7196) );
  AOI22_X1 U4475 ( .A1(reg_mem[295]), .A2(n2660), .B1(n7197), .B2(data_w[7]), 
        .ZN(n2667) );
  INV_X1 U4476 ( .A(n2668), .ZN(n8918) );
  AOI22_X1 U4477 ( .A1(reg_mem[296]), .A2(n2669), .B1(n8926), .B2(data_w[0]), 
        .ZN(n2668) );
  INV_X1 U4478 ( .A(n2670), .ZN(n8919) );
  AOI22_X1 U4479 ( .A1(reg_mem[297]), .A2(n2669), .B1(n8926), .B2(data_w[1]), 
        .ZN(n2670) );
  INV_X1 U4480 ( .A(n2671), .ZN(n8920) );
  AOI22_X1 U4481 ( .A1(reg_mem[298]), .A2(n2669), .B1(n8926), .B2(data_w[2]), 
        .ZN(n2671) );
  INV_X1 U4482 ( .A(n2672), .ZN(n8921) );
  AOI22_X1 U4483 ( .A1(reg_mem[299]), .A2(n2669), .B1(n8926), .B2(data_w[3]), 
        .ZN(n2672) );
  INV_X1 U4484 ( .A(n2673), .ZN(n8922) );
  AOI22_X1 U4485 ( .A1(reg_mem[300]), .A2(n2669), .B1(n8926), .B2(data_w[4]), 
        .ZN(n2673) );
  INV_X1 U4486 ( .A(n2674), .ZN(n8923) );
  AOI22_X1 U4487 ( .A1(reg_mem[301]), .A2(n2669), .B1(n8926), .B2(data_w[5]), 
        .ZN(n2674) );
  INV_X1 U4488 ( .A(n2675), .ZN(n8924) );
  AOI22_X1 U4489 ( .A1(reg_mem[302]), .A2(n2669), .B1(n8926), .B2(data_w[6]), 
        .ZN(n2675) );
  INV_X1 U4490 ( .A(n2676), .ZN(n8925) );
  AOI22_X1 U4491 ( .A1(reg_mem[303]), .A2(n2669), .B1(n8926), .B2(data_w[7]), 
        .ZN(n2676) );
  INV_X1 U4492 ( .A(n2677), .ZN(n7765) );
  AOI22_X1 U4493 ( .A1(reg_mem[304]), .A2(n2678), .B1(n7773), .B2(data_w[0]), 
        .ZN(n2677) );
  INV_X1 U4494 ( .A(n2679), .ZN(n7766) );
  AOI22_X1 U4495 ( .A1(reg_mem[305]), .A2(n2678), .B1(n7773), .B2(data_w[1]), 
        .ZN(n2679) );
  INV_X1 U4496 ( .A(n2680), .ZN(n7767) );
  AOI22_X1 U4497 ( .A1(reg_mem[306]), .A2(n2678), .B1(n7773), .B2(data_w[2]), 
        .ZN(n2680) );
  INV_X1 U4498 ( .A(n2681), .ZN(n7768) );
  AOI22_X1 U4499 ( .A1(reg_mem[307]), .A2(n2678), .B1(n7773), .B2(data_w[3]), 
        .ZN(n2681) );
  INV_X1 U4500 ( .A(n2682), .ZN(n7769) );
  AOI22_X1 U4501 ( .A1(reg_mem[308]), .A2(n2678), .B1(n7773), .B2(data_w[4]), 
        .ZN(n2682) );
  INV_X1 U4502 ( .A(n2683), .ZN(n7770) );
  AOI22_X1 U4503 ( .A1(reg_mem[309]), .A2(n2678), .B1(n7773), .B2(data_w[5]), 
        .ZN(n2683) );
  INV_X1 U4504 ( .A(n2684), .ZN(n7771) );
  AOI22_X1 U4505 ( .A1(reg_mem[310]), .A2(n2678), .B1(n7773), .B2(data_w[6]), 
        .ZN(n2684) );
  INV_X1 U4506 ( .A(n2685), .ZN(n7772) );
  AOI22_X1 U4507 ( .A1(reg_mem[311]), .A2(n2678), .B1(n7773), .B2(data_w[7]), 
        .ZN(n2685) );
  INV_X1 U4508 ( .A(n2686), .ZN(n8342) );
  AOI22_X1 U4509 ( .A1(reg_mem[312]), .A2(n2687), .B1(n8350), .B2(data_w[0]), 
        .ZN(n2686) );
  INV_X1 U4510 ( .A(n2688), .ZN(n8343) );
  AOI22_X1 U4511 ( .A1(reg_mem[313]), .A2(n2687), .B1(n8350), .B2(data_w[1]), 
        .ZN(n2688) );
  INV_X1 U4512 ( .A(n2689), .ZN(n8344) );
  AOI22_X1 U4513 ( .A1(reg_mem[314]), .A2(n2687), .B1(n8350), .B2(data_w[2]), 
        .ZN(n2689) );
  INV_X1 U4514 ( .A(n2690), .ZN(n8345) );
  AOI22_X1 U4515 ( .A1(reg_mem[315]), .A2(n2687), .B1(n8350), .B2(data_w[3]), 
        .ZN(n2690) );
  INV_X1 U4516 ( .A(n2691), .ZN(n8346) );
  AOI22_X1 U4517 ( .A1(reg_mem[316]), .A2(n2687), .B1(n8350), .B2(data_w[4]), 
        .ZN(n2691) );
  INV_X1 U4518 ( .A(n2692), .ZN(n8347) );
  AOI22_X1 U4519 ( .A1(reg_mem[317]), .A2(n2687), .B1(n8350), .B2(data_w[5]), 
        .ZN(n2692) );
  INV_X1 U4520 ( .A(n2693), .ZN(n8348) );
  AOI22_X1 U4521 ( .A1(reg_mem[318]), .A2(n2687), .B1(n8350), .B2(data_w[6]), 
        .ZN(n2693) );
  INV_X1 U4522 ( .A(n2694), .ZN(n8349) );
  AOI22_X1 U4523 ( .A1(reg_mem[319]), .A2(n2687), .B1(n8350), .B2(data_w[7]), 
        .ZN(n2694) );
  INV_X1 U4524 ( .A(n2695), .ZN(n7045) );
  AOI22_X1 U4525 ( .A1(reg_mem[320]), .A2(n2696), .B1(n7053), .B2(data_w[0]), 
        .ZN(n2695) );
  INV_X1 U4526 ( .A(n2697), .ZN(n7046) );
  AOI22_X1 U4527 ( .A1(reg_mem[321]), .A2(n2696), .B1(n7053), .B2(data_w[1]), 
        .ZN(n2697) );
  INV_X1 U4528 ( .A(n2698), .ZN(n7047) );
  AOI22_X1 U4529 ( .A1(reg_mem[322]), .A2(n2696), .B1(n7053), .B2(data_w[2]), 
        .ZN(n2698) );
  INV_X1 U4530 ( .A(n2699), .ZN(n7048) );
  AOI22_X1 U4531 ( .A1(reg_mem[323]), .A2(n2696), .B1(n7053), .B2(data_w[3]), 
        .ZN(n2699) );
  INV_X1 U4532 ( .A(n2700), .ZN(n7049) );
  AOI22_X1 U4533 ( .A1(reg_mem[324]), .A2(n2696), .B1(n7053), .B2(data_w[4]), 
        .ZN(n2700) );
  INV_X1 U4534 ( .A(n2701), .ZN(n7050) );
  AOI22_X1 U4535 ( .A1(reg_mem[325]), .A2(n2696), .B1(n7053), .B2(data_w[5]), 
        .ZN(n2701) );
  INV_X1 U4536 ( .A(n2702), .ZN(n7051) );
  AOI22_X1 U4537 ( .A1(reg_mem[326]), .A2(n2696), .B1(n7053), .B2(data_w[6]), 
        .ZN(n2702) );
  INV_X1 U4538 ( .A(n2703), .ZN(n7052) );
  AOI22_X1 U4539 ( .A1(reg_mem[327]), .A2(n2696), .B1(n7053), .B2(data_w[7]), 
        .ZN(n2703) );
  INV_X1 U4540 ( .A(n2704), .ZN(n8774) );
  AOI22_X1 U4541 ( .A1(reg_mem[328]), .A2(n2705), .B1(n8782), .B2(data_w[0]), 
        .ZN(n2704) );
  INV_X1 U4542 ( .A(n2706), .ZN(n8775) );
  AOI22_X1 U4543 ( .A1(reg_mem[329]), .A2(n2705), .B1(n8782), .B2(data_w[1]), 
        .ZN(n2706) );
  INV_X1 U4544 ( .A(n2707), .ZN(n8776) );
  AOI22_X1 U4545 ( .A1(reg_mem[330]), .A2(n2705), .B1(n8782), .B2(data_w[2]), 
        .ZN(n2707) );
  INV_X1 U4546 ( .A(n2708), .ZN(n8777) );
  AOI22_X1 U4547 ( .A1(reg_mem[331]), .A2(n2705), .B1(n8782), .B2(data_w[3]), 
        .ZN(n2708) );
  INV_X1 U4548 ( .A(n2709), .ZN(n8778) );
  AOI22_X1 U4549 ( .A1(reg_mem[332]), .A2(n2705), .B1(n8782), .B2(data_w[4]), 
        .ZN(n2709) );
  INV_X1 U4550 ( .A(n2710), .ZN(n8779) );
  AOI22_X1 U4551 ( .A1(reg_mem[333]), .A2(n2705), .B1(n8782), .B2(data_w[5]), 
        .ZN(n2710) );
  INV_X1 U4552 ( .A(n2711), .ZN(n8780) );
  AOI22_X1 U4553 ( .A1(reg_mem[334]), .A2(n2705), .B1(n8782), .B2(data_w[6]), 
        .ZN(n2711) );
  INV_X1 U4554 ( .A(n2712), .ZN(n8781) );
  AOI22_X1 U4555 ( .A1(reg_mem[335]), .A2(n2705), .B1(n8782), .B2(data_w[7]), 
        .ZN(n2712) );
  INV_X1 U4556 ( .A(n2713), .ZN(n7621) );
  AOI22_X1 U4557 ( .A1(reg_mem[336]), .A2(n2714), .B1(n7629), .B2(data_w[0]), 
        .ZN(n2713) );
  INV_X1 U4558 ( .A(n2715), .ZN(n7622) );
  AOI22_X1 U4559 ( .A1(reg_mem[337]), .A2(n2714), .B1(n7629), .B2(data_w[1]), 
        .ZN(n2715) );
  INV_X1 U4560 ( .A(n2716), .ZN(n7623) );
  AOI22_X1 U4561 ( .A1(reg_mem[338]), .A2(n2714), .B1(n7629), .B2(data_w[2]), 
        .ZN(n2716) );
  INV_X1 U4562 ( .A(n2717), .ZN(n7624) );
  AOI22_X1 U4563 ( .A1(reg_mem[339]), .A2(n2714), .B1(n7629), .B2(data_w[3]), 
        .ZN(n2717) );
  INV_X1 U4564 ( .A(n2718), .ZN(n7625) );
  AOI22_X1 U4565 ( .A1(reg_mem[340]), .A2(n2714), .B1(n7629), .B2(data_w[4]), 
        .ZN(n2718) );
  INV_X1 U4566 ( .A(n2719), .ZN(n7626) );
  AOI22_X1 U4567 ( .A1(reg_mem[341]), .A2(n2714), .B1(n7629), .B2(data_w[5]), 
        .ZN(n2719) );
  INV_X1 U4568 ( .A(n2720), .ZN(n7627) );
  AOI22_X1 U4569 ( .A1(reg_mem[342]), .A2(n2714), .B1(n7629), .B2(data_w[6]), 
        .ZN(n2720) );
  INV_X1 U4570 ( .A(n2721), .ZN(n7628) );
  AOI22_X1 U4571 ( .A1(reg_mem[343]), .A2(n2714), .B1(n7629), .B2(data_w[7]), 
        .ZN(n2721) );
  INV_X1 U4572 ( .A(n2722), .ZN(n8198) );
  AOI22_X1 U4573 ( .A1(reg_mem[344]), .A2(n2723), .B1(n8206), .B2(data_w[0]), 
        .ZN(n2722) );
  INV_X1 U4574 ( .A(n2724), .ZN(n8199) );
  AOI22_X1 U4575 ( .A1(reg_mem[345]), .A2(n2723), .B1(n8206), .B2(data_w[1]), 
        .ZN(n2724) );
  INV_X1 U4576 ( .A(n2725), .ZN(n8200) );
  AOI22_X1 U4577 ( .A1(reg_mem[346]), .A2(n2723), .B1(n8206), .B2(data_w[2]), 
        .ZN(n2725) );
  INV_X1 U4578 ( .A(n2726), .ZN(n8201) );
  AOI22_X1 U4579 ( .A1(reg_mem[347]), .A2(n2723), .B1(n8206), .B2(data_w[3]), 
        .ZN(n2726) );
  INV_X1 U4580 ( .A(n2727), .ZN(n8202) );
  AOI22_X1 U4581 ( .A1(reg_mem[348]), .A2(n2723), .B1(n8206), .B2(data_w[4]), 
        .ZN(n2727) );
  INV_X1 U4582 ( .A(n2728), .ZN(n8203) );
  AOI22_X1 U4583 ( .A1(reg_mem[349]), .A2(n2723), .B1(n8206), .B2(data_w[5]), 
        .ZN(n2728) );
  INV_X1 U4584 ( .A(n2729), .ZN(n8204) );
  AOI22_X1 U4585 ( .A1(reg_mem[350]), .A2(n2723), .B1(n8206), .B2(data_w[6]), 
        .ZN(n2729) );
  INV_X1 U4586 ( .A(n2730), .ZN(n8205) );
  AOI22_X1 U4587 ( .A1(reg_mem[351]), .A2(n2723), .B1(n8206), .B2(data_w[7]), 
        .ZN(n2730) );
  INV_X1 U4588 ( .A(n2731), .ZN(n6901) );
  AOI22_X1 U4589 ( .A1(reg_mem[352]), .A2(n2732), .B1(n6909), .B2(data_w[0]), 
        .ZN(n2731) );
  INV_X1 U4590 ( .A(n2733), .ZN(n6902) );
  AOI22_X1 U4591 ( .A1(reg_mem[353]), .A2(n2732), .B1(n6909), .B2(data_w[1]), 
        .ZN(n2733) );
  INV_X1 U4592 ( .A(n2734), .ZN(n6903) );
  AOI22_X1 U4593 ( .A1(reg_mem[354]), .A2(n2732), .B1(n6909), .B2(data_w[2]), 
        .ZN(n2734) );
  INV_X1 U4594 ( .A(n2735), .ZN(n6904) );
  AOI22_X1 U4595 ( .A1(reg_mem[355]), .A2(n2732), .B1(n6909), .B2(data_w[3]), 
        .ZN(n2735) );
  INV_X1 U4596 ( .A(n2736), .ZN(n6905) );
  AOI22_X1 U4597 ( .A1(reg_mem[356]), .A2(n2732), .B1(n6909), .B2(data_w[4]), 
        .ZN(n2736) );
  INV_X1 U4598 ( .A(n2737), .ZN(n6906) );
  AOI22_X1 U4599 ( .A1(reg_mem[357]), .A2(n2732), .B1(n6909), .B2(data_w[5]), 
        .ZN(n2737) );
  INV_X1 U4600 ( .A(n2738), .ZN(n6907) );
  AOI22_X1 U4601 ( .A1(reg_mem[358]), .A2(n2732), .B1(n6909), .B2(data_w[6]), 
        .ZN(n2738) );
  INV_X1 U4602 ( .A(n2739), .ZN(n6908) );
  AOI22_X1 U4603 ( .A1(reg_mem[359]), .A2(n2732), .B1(n6909), .B2(data_w[7]), 
        .ZN(n2739) );
  INV_X1 U4604 ( .A(n2740), .ZN(n8630) );
  AOI22_X1 U4605 ( .A1(reg_mem[360]), .A2(n2741), .B1(n8638), .B2(data_w[0]), 
        .ZN(n2740) );
  INV_X1 U4606 ( .A(n2742), .ZN(n8631) );
  AOI22_X1 U4607 ( .A1(reg_mem[361]), .A2(n2741), .B1(n8638), .B2(data_w[1]), 
        .ZN(n2742) );
  INV_X1 U4608 ( .A(n2743), .ZN(n8632) );
  AOI22_X1 U4609 ( .A1(reg_mem[362]), .A2(n2741), .B1(n8638), .B2(data_w[2]), 
        .ZN(n2743) );
  INV_X1 U4610 ( .A(n2744), .ZN(n8633) );
  AOI22_X1 U4611 ( .A1(reg_mem[363]), .A2(n2741), .B1(n8638), .B2(data_w[3]), 
        .ZN(n2744) );
  INV_X1 U4612 ( .A(n2745), .ZN(n8634) );
  AOI22_X1 U4613 ( .A1(reg_mem[364]), .A2(n2741), .B1(n8638), .B2(data_w[4]), 
        .ZN(n2745) );
  INV_X1 U4614 ( .A(n2746), .ZN(n8635) );
  AOI22_X1 U4615 ( .A1(reg_mem[365]), .A2(n2741), .B1(n8638), .B2(data_w[5]), 
        .ZN(n2746) );
  INV_X1 U4616 ( .A(n2747), .ZN(n8636) );
  AOI22_X1 U4617 ( .A1(reg_mem[366]), .A2(n2741), .B1(n8638), .B2(data_w[6]), 
        .ZN(n2747) );
  INV_X1 U4618 ( .A(n2748), .ZN(n8637) );
  AOI22_X1 U4619 ( .A1(reg_mem[367]), .A2(n2741), .B1(n8638), .B2(data_w[7]), 
        .ZN(n2748) );
  INV_X1 U4620 ( .A(n2749), .ZN(n7477) );
  AOI22_X1 U4621 ( .A1(reg_mem[368]), .A2(n2750), .B1(n7485), .B2(data_w[0]), 
        .ZN(n2749) );
  INV_X1 U4622 ( .A(n2751), .ZN(n7478) );
  AOI22_X1 U4623 ( .A1(reg_mem[369]), .A2(n2750), .B1(n7485), .B2(data_w[1]), 
        .ZN(n2751) );
  INV_X1 U4624 ( .A(n2752), .ZN(n7479) );
  AOI22_X1 U4625 ( .A1(reg_mem[370]), .A2(n2750), .B1(n7485), .B2(data_w[2]), 
        .ZN(n2752) );
  INV_X1 U4626 ( .A(n2753), .ZN(n7480) );
  AOI22_X1 U4627 ( .A1(reg_mem[371]), .A2(n2750), .B1(n7485), .B2(data_w[3]), 
        .ZN(n2753) );
  INV_X1 U4628 ( .A(n2754), .ZN(n7481) );
  AOI22_X1 U4629 ( .A1(reg_mem[372]), .A2(n2750), .B1(n7485), .B2(data_w[4]), 
        .ZN(n2754) );
  INV_X1 U4630 ( .A(n2755), .ZN(n7482) );
  AOI22_X1 U4631 ( .A1(reg_mem[373]), .A2(n2750), .B1(n7485), .B2(data_w[5]), 
        .ZN(n2755) );
  INV_X1 U4632 ( .A(n2756), .ZN(n7483) );
  AOI22_X1 U4633 ( .A1(reg_mem[374]), .A2(n2750), .B1(n7485), .B2(data_w[6]), 
        .ZN(n2756) );
  INV_X1 U4634 ( .A(n2757), .ZN(n7484) );
  AOI22_X1 U4635 ( .A1(reg_mem[375]), .A2(n2750), .B1(n7485), .B2(data_w[7]), 
        .ZN(n2757) );
  INV_X1 U4636 ( .A(n2758), .ZN(n8054) );
  AOI22_X1 U4637 ( .A1(reg_mem[376]), .A2(n2759), .B1(n8062), .B2(data_w[0]), 
        .ZN(n2758) );
  INV_X1 U4638 ( .A(n2760), .ZN(n8055) );
  AOI22_X1 U4639 ( .A1(reg_mem[377]), .A2(n2759), .B1(n8062), .B2(data_w[1]), 
        .ZN(n2760) );
  INV_X1 U4640 ( .A(n2761), .ZN(n8056) );
  AOI22_X1 U4641 ( .A1(reg_mem[378]), .A2(n2759), .B1(n8062), .B2(data_w[2]), 
        .ZN(n2761) );
  INV_X1 U4642 ( .A(n2762), .ZN(n8057) );
  AOI22_X1 U4643 ( .A1(reg_mem[379]), .A2(n2759), .B1(n8062), .B2(data_w[3]), 
        .ZN(n2762) );
  INV_X1 U4644 ( .A(n2763), .ZN(n8058) );
  AOI22_X1 U4645 ( .A1(reg_mem[380]), .A2(n2759), .B1(n8062), .B2(data_w[4]), 
        .ZN(n2763) );
  INV_X1 U4646 ( .A(n2764), .ZN(n8059) );
  AOI22_X1 U4647 ( .A1(reg_mem[381]), .A2(n2759), .B1(n8062), .B2(data_w[5]), 
        .ZN(n2764) );
  INV_X1 U4648 ( .A(n2765), .ZN(n8060) );
  AOI22_X1 U4649 ( .A1(reg_mem[382]), .A2(n2759), .B1(n8062), .B2(data_w[6]), 
        .ZN(n2765) );
  INV_X1 U4650 ( .A(n2766), .ZN(n8061) );
  AOI22_X1 U4651 ( .A1(reg_mem[383]), .A2(n2759), .B1(n8062), .B2(data_w[7]), 
        .ZN(n2766) );
  INV_X1 U4652 ( .A(n2768), .ZN(n7324) );
  AOI22_X1 U4653 ( .A1(reg_mem[384]), .A2(n2769), .B1(n7332), .B2(data_w[0]), 
        .ZN(n2768) );
  INV_X1 U4654 ( .A(n2770), .ZN(n7325) );
  AOI22_X1 U4655 ( .A1(reg_mem[385]), .A2(n2769), .B1(n7332), .B2(data_w[1]), 
        .ZN(n2770) );
  INV_X1 U4656 ( .A(n2771), .ZN(n7326) );
  AOI22_X1 U4657 ( .A1(reg_mem[386]), .A2(n2769), .B1(n7332), .B2(data_w[2]), 
        .ZN(n2771) );
  INV_X1 U4658 ( .A(n2772), .ZN(n7327) );
  AOI22_X1 U4659 ( .A1(reg_mem[387]), .A2(n2769), .B1(n7332), .B2(data_w[3]), 
        .ZN(n2772) );
  INV_X1 U4660 ( .A(n2773), .ZN(n7328) );
  AOI22_X1 U4661 ( .A1(reg_mem[388]), .A2(n2769), .B1(n7332), .B2(data_w[4]), 
        .ZN(n2773) );
  INV_X1 U4662 ( .A(n2774), .ZN(n7329) );
  AOI22_X1 U4663 ( .A1(reg_mem[389]), .A2(n2769), .B1(n7332), .B2(data_w[5]), 
        .ZN(n2774) );
  INV_X1 U4664 ( .A(n2775), .ZN(n7330) );
  AOI22_X1 U4665 ( .A1(reg_mem[390]), .A2(n2769), .B1(n7332), .B2(data_w[6]), 
        .ZN(n2775) );
  INV_X1 U4666 ( .A(n2776), .ZN(n7331) );
  AOI22_X1 U4667 ( .A1(reg_mem[391]), .A2(n2769), .B1(n7332), .B2(data_w[7]), 
        .ZN(n2776) );
  INV_X1 U4668 ( .A(n2778), .ZN(n9053) );
  AOI22_X1 U4669 ( .A1(reg_mem[392]), .A2(n2779), .B1(n9061), .B2(data_w[0]), 
        .ZN(n2778) );
  INV_X1 U4670 ( .A(n2780), .ZN(n9054) );
  AOI22_X1 U4671 ( .A1(reg_mem[393]), .A2(n2779), .B1(n9061), .B2(data_w[1]), 
        .ZN(n2780) );
  INV_X1 U4672 ( .A(n2781), .ZN(n9055) );
  AOI22_X1 U4673 ( .A1(reg_mem[394]), .A2(n2779), .B1(n9061), .B2(data_w[2]), 
        .ZN(n2781) );
  INV_X1 U4674 ( .A(n2782), .ZN(n9056) );
  AOI22_X1 U4675 ( .A1(reg_mem[395]), .A2(n2779), .B1(n9061), .B2(data_w[3]), 
        .ZN(n2782) );
  INV_X1 U4676 ( .A(n2783), .ZN(n9057) );
  AOI22_X1 U4677 ( .A1(reg_mem[396]), .A2(n2779), .B1(n9061), .B2(data_w[4]), 
        .ZN(n2783) );
  INV_X1 U4678 ( .A(n2784), .ZN(n9058) );
  AOI22_X1 U4679 ( .A1(reg_mem[397]), .A2(n2779), .B1(n9061), .B2(data_w[5]), 
        .ZN(n2784) );
  INV_X1 U4680 ( .A(n2785), .ZN(n9059) );
  AOI22_X1 U4681 ( .A1(reg_mem[398]), .A2(n2779), .B1(n9061), .B2(data_w[6]), 
        .ZN(n2785) );
  INV_X1 U4682 ( .A(n2786), .ZN(n9060) );
  AOI22_X1 U4683 ( .A1(reg_mem[399]), .A2(n2779), .B1(n9061), .B2(data_w[7]), 
        .ZN(n2786) );
  INV_X1 U4684 ( .A(n2787), .ZN(n7900) );
  AOI22_X1 U4685 ( .A1(reg_mem[400]), .A2(n2788), .B1(n7908), .B2(data_w[0]), 
        .ZN(n2787) );
  INV_X1 U4686 ( .A(n2789), .ZN(n7901) );
  AOI22_X1 U4687 ( .A1(reg_mem[401]), .A2(n2788), .B1(n7908), .B2(data_w[1]), 
        .ZN(n2789) );
  INV_X1 U4688 ( .A(n2790), .ZN(n7902) );
  AOI22_X1 U4689 ( .A1(reg_mem[402]), .A2(n2788), .B1(n7908), .B2(data_w[2]), 
        .ZN(n2790) );
  INV_X1 U4690 ( .A(n2791), .ZN(n7903) );
  AOI22_X1 U4691 ( .A1(reg_mem[403]), .A2(n2788), .B1(n7908), .B2(data_w[3]), 
        .ZN(n2791) );
  INV_X1 U4692 ( .A(n2792), .ZN(n7904) );
  AOI22_X1 U4693 ( .A1(reg_mem[404]), .A2(n2788), .B1(n7908), .B2(data_w[4]), 
        .ZN(n2792) );
  INV_X1 U4694 ( .A(n2793), .ZN(n7905) );
  AOI22_X1 U4695 ( .A1(reg_mem[405]), .A2(n2788), .B1(n7908), .B2(data_w[5]), 
        .ZN(n2793) );
  INV_X1 U4696 ( .A(n2794), .ZN(n7906) );
  AOI22_X1 U4697 ( .A1(reg_mem[406]), .A2(n2788), .B1(n7908), .B2(data_w[6]), 
        .ZN(n2794) );
  INV_X1 U4698 ( .A(n2795), .ZN(n7907) );
  AOI22_X1 U4699 ( .A1(reg_mem[407]), .A2(n2788), .B1(n7908), .B2(data_w[7]), 
        .ZN(n2795) );
  INV_X1 U4700 ( .A(n2796), .ZN(n8477) );
  AOI22_X1 U4701 ( .A1(reg_mem[408]), .A2(n2797), .B1(n8485), .B2(data_w[0]), 
        .ZN(n2796) );
  INV_X1 U4702 ( .A(n2798), .ZN(n8478) );
  AOI22_X1 U4703 ( .A1(reg_mem[409]), .A2(n2797), .B1(n8485), .B2(data_w[1]), 
        .ZN(n2798) );
  INV_X1 U4704 ( .A(n2799), .ZN(n8479) );
  AOI22_X1 U4705 ( .A1(reg_mem[410]), .A2(n2797), .B1(n8485), .B2(data_w[2]), 
        .ZN(n2799) );
  INV_X1 U4706 ( .A(n2800), .ZN(n8480) );
  AOI22_X1 U4707 ( .A1(reg_mem[411]), .A2(n2797), .B1(n8485), .B2(data_w[3]), 
        .ZN(n2800) );
  INV_X1 U4708 ( .A(n2801), .ZN(n8481) );
  AOI22_X1 U4709 ( .A1(reg_mem[412]), .A2(n2797), .B1(n8485), .B2(data_w[4]), 
        .ZN(n2801) );
  INV_X1 U4710 ( .A(n2802), .ZN(n8482) );
  AOI22_X1 U4711 ( .A1(reg_mem[413]), .A2(n2797), .B1(n8485), .B2(data_w[5]), 
        .ZN(n2802) );
  INV_X1 U4712 ( .A(n2803), .ZN(n8483) );
  AOI22_X1 U4713 ( .A1(reg_mem[414]), .A2(n2797), .B1(n8485), .B2(data_w[6]), 
        .ZN(n2803) );
  INV_X1 U4714 ( .A(n2804), .ZN(n8484) );
  AOI22_X1 U4715 ( .A1(reg_mem[415]), .A2(n2797), .B1(n8485), .B2(data_w[7]), 
        .ZN(n2804) );
  MUX2_X1 U4716 ( .A(reg_mem[8]), .B(reg_mem[0]), .S(n6762), .Z(n4665) );
  MUX2_X1 U4717 ( .A(reg_mem[24]), .B(reg_mem[16]), .S(n6779), .Z(n4666) );
  MUX2_X1 U4718 ( .A(n4666), .B(n4665), .S(n6722), .Z(n4667) );
  MUX2_X1 U4719 ( .A(reg_mem[40]), .B(reg_mem[32]), .S(n6753), .Z(n4668) );
  MUX2_X1 U4720 ( .A(reg_mem[56]), .B(reg_mem[48]), .S(n6745), .Z(n4669) );
  MUX2_X1 U4721 ( .A(n4669), .B(n4668), .S(n6724), .Z(n4670) );
  MUX2_X1 U4722 ( .A(n4670), .B(n4667), .S(n6707), .Z(n4671) );
  MUX2_X1 U4723 ( .A(reg_mem[72]), .B(reg_mem[64]), .S(n6762), .Z(n4672) );
  MUX2_X1 U4724 ( .A(reg_mem[88]), .B(reg_mem[80]), .S(n6778), .Z(n4673) );
  MUX2_X1 U4725 ( .A(n4673), .B(n4672), .S(n6723), .Z(n4674) );
  MUX2_X1 U4726 ( .A(reg_mem[104]), .B(reg_mem[96]), .S(n6740), .Z(n4675) );
  MUX2_X1 U4727 ( .A(reg_mem[120]), .B(reg_mem[112]), .S(n6741), .Z(n4676) );
  MUX2_X1 U4728 ( .A(n4676), .B(n4675), .S(n6723), .Z(n4677) );
  MUX2_X1 U4729 ( .A(n4677), .B(n4674), .S(n6717), .Z(n4678) );
  MUX2_X1 U4730 ( .A(n4678), .B(n4671), .S(n6704), .Z(n4679) );
  MUX2_X1 U4731 ( .A(reg_mem[136]), .B(reg_mem[128]), .S(n6741), .Z(n4680) );
  MUX2_X1 U4732 ( .A(reg_mem[152]), .B(reg_mem[144]), .S(n6773), .Z(n4681) );
  MUX2_X1 U4733 ( .A(n4681), .B(n4680), .S(n6723), .Z(n4682) );
  MUX2_X1 U4734 ( .A(reg_mem[168]), .B(reg_mem[160]), .S(n6740), .Z(n4683) );
  MUX2_X1 U4735 ( .A(reg_mem[184]), .B(reg_mem[176]), .S(n6741), .Z(n4684) );
  MUX2_X1 U4736 ( .A(n4684), .B(n4683), .S(n6722), .Z(n4685) );
  MUX2_X1 U4737 ( .A(n4685), .B(n4682), .S(addr_r[2]), .Z(n4686) );
  MUX2_X1 U4738 ( .A(reg_mem[200]), .B(reg_mem[192]), .S(n6760), .Z(n4687) );
  MUX2_X1 U4739 ( .A(reg_mem[216]), .B(reg_mem[208]), .S(n6781), .Z(n4688) );
  MUX2_X1 U4740 ( .A(n4688), .B(n4687), .S(n6724), .Z(n4689) );
  MUX2_X1 U4741 ( .A(reg_mem[232]), .B(reg_mem[224]), .S(n6780), .Z(n4690) );
  MUX2_X1 U4742 ( .A(reg_mem[248]), .B(reg_mem[240]), .S(n6759), .Z(n4691) );
  MUX2_X1 U4743 ( .A(n4691), .B(n4690), .S(n6722), .Z(n4692) );
  MUX2_X1 U4744 ( .A(n4692), .B(n4689), .S(n6709), .Z(n4693) );
  MUX2_X1 U4745 ( .A(n4693), .B(n4686), .S(n6701), .Z(n4694) );
  MUX2_X1 U4746 ( .A(n4694), .B(n4679), .S(n6699), .Z(n4695) );
  MUX2_X1 U4747 ( .A(reg_mem[264]), .B(reg_mem[256]), .S(n6742), .Z(n4696) );
  MUX2_X1 U4748 ( .A(reg_mem[280]), .B(reg_mem[272]), .S(n6741), .Z(n4697) );
  MUX2_X1 U4749 ( .A(n4697), .B(n4696), .S(n6721), .Z(n4698) );
  MUX2_X1 U4750 ( .A(reg_mem[296]), .B(reg_mem[288]), .S(n6755), .Z(n4699) );
  MUX2_X1 U4751 ( .A(reg_mem[312]), .B(reg_mem[304]), .S(n6773), .Z(n4700) );
  MUX2_X1 U4752 ( .A(n4700), .B(n4699), .S(n6725), .Z(n4701) );
  MUX2_X1 U4753 ( .A(n4701), .B(n4698), .S(n6711), .Z(n4702) );
  MUX2_X1 U4754 ( .A(reg_mem[328]), .B(reg_mem[320]), .S(n6769), .Z(n4703) );
  MUX2_X1 U4755 ( .A(reg_mem[344]), .B(reg_mem[336]), .S(n6742), .Z(n4704) );
  MUX2_X1 U4756 ( .A(n4704), .B(n4703), .S(n6723), .Z(n4705) );
  MUX2_X1 U4757 ( .A(reg_mem[360]), .B(reg_mem[352]), .S(n6774), .Z(n4706) );
  MUX2_X1 U4758 ( .A(reg_mem[376]), .B(reg_mem[368]), .S(n6760), .Z(n4707) );
  MUX2_X1 U4759 ( .A(n4707), .B(n4706), .S(n6725), .Z(n4708) );
  MUX2_X1 U4760 ( .A(n4708), .B(n4705), .S(n6711), .Z(n4709) );
  MUX2_X1 U4761 ( .A(n4709), .B(n4702), .S(n6705), .Z(n4710) );
  MUX2_X1 U4762 ( .A(reg_mem[392]), .B(reg_mem[384]), .S(n6756), .Z(n4711) );
  MUX2_X1 U4763 ( .A(reg_mem[408]), .B(reg_mem[400]), .S(n6761), .Z(n4712) );
  MUX2_X1 U4764 ( .A(n4712), .B(n4711), .S(n6721), .Z(n4713) );
  MUX2_X1 U4765 ( .A(reg_mem[424]), .B(reg_mem[416]), .S(n6783), .Z(n4714) );
  MUX2_X1 U4766 ( .A(reg_mem[440]), .B(reg_mem[432]), .S(n6779), .Z(n4715) );
  MUX2_X1 U4767 ( .A(n4715), .B(n4714), .S(n6718), .Z(n4716) );
  MUX2_X1 U4768 ( .A(n4716), .B(n4713), .S(n6716), .Z(n4717) );
  MUX2_X1 U4769 ( .A(reg_mem[456]), .B(reg_mem[448]), .S(n6740), .Z(n4718) );
  MUX2_X1 U4770 ( .A(reg_mem[472]), .B(reg_mem[464]), .S(n6768), .Z(n4719) );
  MUX2_X1 U4771 ( .A(n4719), .B(n4718), .S(n6721), .Z(n4720) );
  MUX2_X1 U4772 ( .A(reg_mem[488]), .B(reg_mem[480]), .S(n6783), .Z(n4721) );
  MUX2_X1 U4773 ( .A(reg_mem[504]), .B(reg_mem[496]), .S(n6760), .Z(n4722) );
  MUX2_X1 U4774 ( .A(n4722), .B(n4721), .S(n6735), .Z(n4723) );
  MUX2_X1 U4775 ( .A(n4723), .B(n4720), .S(n6713), .Z(n4724) );
  MUX2_X1 U4776 ( .A(n4724), .B(n4717), .S(n6703), .Z(n4725) );
  MUX2_X1 U4777 ( .A(n4725), .B(n4710), .S(n6699), .Z(n4726) );
  MUX2_X1 U4778 ( .A(n4726), .B(n4695), .S(n6697), .Z(n4727) );
  MUX2_X1 U4779 ( .A(reg_mem[520]), .B(reg_mem[512]), .S(n6783), .Z(n4728) );
  MUX2_X1 U4780 ( .A(reg_mem[536]), .B(reg_mem[528]), .S(n6740), .Z(n4729) );
  MUX2_X1 U4781 ( .A(n4729), .B(n4728), .S(n6734), .Z(n4730) );
  MUX2_X1 U4782 ( .A(reg_mem[552]), .B(reg_mem[544]), .S(n6744), .Z(n4731) );
  MUX2_X1 U4783 ( .A(reg_mem[568]), .B(reg_mem[560]), .S(n6783), .Z(n4732) );
  MUX2_X1 U4784 ( .A(n4732), .B(n4731), .S(n6721), .Z(n4733) );
  MUX2_X1 U4785 ( .A(n4733), .B(n4730), .S(n6715), .Z(n4734) );
  MUX2_X1 U4786 ( .A(reg_mem[584]), .B(reg_mem[576]), .S(n6763), .Z(n4735) );
  MUX2_X1 U4787 ( .A(reg_mem[600]), .B(reg_mem[592]), .S(n6740), .Z(n4736) );
  MUX2_X1 U4788 ( .A(n4736), .B(n4735), .S(n6720), .Z(n4737) );
  MUX2_X1 U4789 ( .A(reg_mem[616]), .B(reg_mem[608]), .S(n6782), .Z(n4738) );
  MUX2_X1 U4790 ( .A(reg_mem[632]), .B(reg_mem[624]), .S(n6757), .Z(n4739) );
  MUX2_X1 U4791 ( .A(n4739), .B(n4738), .S(n6719), .Z(n4740) );
  MUX2_X1 U4792 ( .A(n4740), .B(n4737), .S(n6714), .Z(n4741) );
  MUX2_X1 U4793 ( .A(n4741), .B(n4734), .S(n6704), .Z(n4742) );
  MUX2_X1 U4794 ( .A(reg_mem[648]), .B(reg_mem[640]), .S(n6740), .Z(n4743) );
  MUX2_X1 U4795 ( .A(reg_mem[664]), .B(reg_mem[656]), .S(n6766), .Z(n4744) );
  MUX2_X1 U4796 ( .A(n4744), .B(n4743), .S(n6735), .Z(n4745) );
  MUX2_X1 U4797 ( .A(reg_mem[680]), .B(reg_mem[672]), .S(n6742), .Z(n4746) );
  MUX2_X1 U4798 ( .A(reg_mem[696]), .B(reg_mem[688]), .S(n6765), .Z(n4747) );
  MUX2_X1 U4799 ( .A(n4747), .B(n4746), .S(n6729), .Z(n4748) );
  MUX2_X1 U4800 ( .A(n4748), .B(n4745), .S(n6713), .Z(n4749) );
  MUX2_X1 U4801 ( .A(reg_mem[712]), .B(reg_mem[704]), .S(n6742), .Z(n4750) );
  MUX2_X1 U4802 ( .A(reg_mem[728]), .B(reg_mem[720]), .S(n6777), .Z(n4751) );
  MUX2_X1 U4803 ( .A(n4751), .B(n4750), .S(n6718), .Z(n4752) );
  MUX2_X1 U4804 ( .A(reg_mem[744]), .B(reg_mem[736]), .S(n6782), .Z(n4753) );
  MUX2_X1 U4805 ( .A(reg_mem[760]), .B(reg_mem[752]), .S(n6770), .Z(n4754) );
  MUX2_X1 U4806 ( .A(n4754), .B(n4753), .S(n6718), .Z(n4755) );
  MUX2_X1 U4807 ( .A(n4755), .B(n4752), .S(addr_r[2]), .Z(n4756) );
  MUX2_X1 U4808 ( .A(n4756), .B(n4749), .S(n6702), .Z(n4757) );
  MUX2_X1 U4809 ( .A(n4757), .B(n4742), .S(addr_r[4]), .Z(n4758) );
  MUX2_X1 U4810 ( .A(reg_mem[776]), .B(reg_mem[768]), .S(n6778), .Z(n4759) );
  MUX2_X1 U4811 ( .A(reg_mem[792]), .B(reg_mem[784]), .S(n6783), .Z(n4760) );
  MUX2_X1 U4812 ( .A(n4760), .B(n4759), .S(n6721), .Z(n4761) );
  MUX2_X1 U4813 ( .A(reg_mem[808]), .B(reg_mem[800]), .S(n6760), .Z(n4762) );
  MUX2_X1 U4814 ( .A(reg_mem[824]), .B(reg_mem[816]), .S(n6772), .Z(n4763) );
  MUX2_X1 U4815 ( .A(n4763), .B(n4762), .S(n6732), .Z(n4764) );
  MUX2_X1 U4816 ( .A(n4764), .B(n4761), .S(n6715), .Z(n4765) );
  MUX2_X1 U4817 ( .A(reg_mem[840]), .B(reg_mem[832]), .S(addr_r[0]), .Z(n4766)
         );
  MUX2_X1 U4818 ( .A(reg_mem[856]), .B(reg_mem[848]), .S(n6783), .Z(n4767) );
  MUX2_X1 U4819 ( .A(n4767), .B(n4766), .S(n6738), .Z(n4768) );
  MUX2_X1 U4820 ( .A(reg_mem[872]), .B(reg_mem[864]), .S(n6779), .Z(n4769) );
  MUX2_X1 U4821 ( .A(reg_mem[888]), .B(reg_mem[880]), .S(addr_r[0]), .Z(n4770)
         );
  MUX2_X1 U4822 ( .A(n4770), .B(n4769), .S(n6734), .Z(n4771) );
  MUX2_X1 U4823 ( .A(n4771), .B(n4768), .S(addr_r[2]), .Z(n4772) );
  MUX2_X1 U4824 ( .A(n4772), .B(n4765), .S(n6705), .Z(n4773) );
  MUX2_X1 U4825 ( .A(reg_mem[904]), .B(reg_mem[896]), .S(n6754), .Z(n4774) );
  MUX2_X1 U4826 ( .A(reg_mem[920]), .B(reg_mem[912]), .S(n6783), .Z(n4775) );
  MUX2_X1 U4827 ( .A(n4775), .B(n4774), .S(n6733), .Z(n4776) );
  MUX2_X1 U4828 ( .A(reg_mem[936]), .B(reg_mem[928]), .S(n6780), .Z(n4777) );
  MUX2_X1 U4829 ( .A(reg_mem[952]), .B(reg_mem[944]), .S(n6775), .Z(n4778) );
  MUX2_X1 U4830 ( .A(n4778), .B(n4777), .S(n6731), .Z(n4779) );
  MUX2_X1 U4831 ( .A(n4779), .B(n4776), .S(n6714), .Z(n4780) );
  MUX2_X1 U4832 ( .A(reg_mem[968]), .B(reg_mem[960]), .S(n6746), .Z(n4781) );
  MUX2_X1 U4833 ( .A(reg_mem[984]), .B(reg_mem[976]), .S(addr_r[0]), .Z(n4782)
         );
  MUX2_X1 U4834 ( .A(n4782), .B(n4781), .S(n6718), .Z(n4783) );
  MUX2_X1 U4835 ( .A(reg_mem[1000]), .B(reg_mem[992]), .S(addr_r[0]), .Z(n4784) );
  MUX2_X1 U4836 ( .A(reg_mem[1016]), .B(reg_mem[1008]), .S(n6781), .Z(n4785)
         );
  MUX2_X1 U4837 ( .A(n4785), .B(n4784), .S(n6733), .Z(n4786) );
  MUX2_X1 U4838 ( .A(n4786), .B(n4783), .S(addr_r[2]), .Z(n4787) );
  MUX2_X1 U4839 ( .A(n4787), .B(n4780), .S(n6706), .Z(n4788) );
  MUX2_X1 U4840 ( .A(n4788), .B(n4773), .S(addr_r[4]), .Z(n4789) );
  MUX2_X1 U4841 ( .A(n4789), .B(n4758), .S(addr_r[5]), .Z(n4790) );
  MUX2_X1 U4842 ( .A(n4790), .B(n4727), .S(addr_r[6]), .Z(n4791) );
  MUX2_X1 U4843 ( .A(reg_mem[1032]), .B(reg_mem[1024]), .S(n6744), .Z(n4792)
         );
  MUX2_X1 U4844 ( .A(reg_mem[1048]), .B(reg_mem[1040]), .S(n6764), .Z(n4793)
         );
  MUX2_X1 U4845 ( .A(n4793), .B(n4792), .S(n6737), .Z(n4794) );
  MUX2_X1 U4846 ( .A(reg_mem[1064]), .B(reg_mem[1056]), .S(n6775), .Z(n4795)
         );
  MUX2_X1 U4847 ( .A(reg_mem[1080]), .B(reg_mem[1072]), .S(n6769), .Z(n4796)
         );
  MUX2_X1 U4848 ( .A(n4796), .B(n4795), .S(n6733), .Z(n4797) );
  MUX2_X1 U4849 ( .A(n4797), .B(n4794), .S(n6708), .Z(n4798) );
  MUX2_X1 U4850 ( .A(reg_mem[1096]), .B(reg_mem[1088]), .S(n6768), .Z(n4799)
         );
  MUX2_X1 U4851 ( .A(reg_mem[1112]), .B(reg_mem[1104]), .S(n6741), .Z(n4800)
         );
  MUX2_X1 U4852 ( .A(n4800), .B(n4799), .S(n6718), .Z(n4801) );
  MUX2_X1 U4853 ( .A(reg_mem[1128]), .B(reg_mem[1120]), .S(n6741), .Z(n4802)
         );
  MUX2_X1 U4854 ( .A(reg_mem[1144]), .B(reg_mem[1136]), .S(n6781), .Z(n4803)
         );
  MUX2_X1 U4855 ( .A(n4803), .B(n4802), .S(n6734), .Z(n4804) );
  MUX2_X1 U4856 ( .A(n4804), .B(n4801), .S(n6707), .Z(n4805) );
  MUX2_X1 U4857 ( .A(n4805), .B(n4798), .S(n6705), .Z(n4806) );
  MUX2_X1 U4858 ( .A(reg_mem[1160]), .B(reg_mem[1152]), .S(n6753), .Z(n4807)
         );
  MUX2_X1 U4859 ( .A(reg_mem[1176]), .B(reg_mem[1168]), .S(n6745), .Z(n4808)
         );
  MUX2_X1 U4860 ( .A(n4808), .B(n4807), .S(n6732), .Z(n4809) );
  MUX2_X1 U4861 ( .A(reg_mem[1192]), .B(reg_mem[1184]), .S(n6755), .Z(n4810)
         );
  MUX2_X1 U4862 ( .A(reg_mem[1208]), .B(reg_mem[1200]), .S(n6740), .Z(n4811)
         );
  MUX2_X1 U4863 ( .A(n4811), .B(n4810), .S(n6735), .Z(n4812) );
  MUX2_X1 U4864 ( .A(n4812), .B(n4809), .S(n6712), .Z(n4813) );
  MUX2_X1 U4865 ( .A(reg_mem[1224]), .B(reg_mem[1216]), .S(n6768), .Z(n4814)
         );
  MUX2_X1 U4866 ( .A(reg_mem[1240]), .B(reg_mem[1232]), .S(n6764), .Z(n4815)
         );
  MUX2_X1 U4867 ( .A(n4815), .B(n4814), .S(n6731), .Z(n4816) );
  MUX2_X1 U4868 ( .A(reg_mem[1256]), .B(reg_mem[1248]), .S(n6772), .Z(n4817)
         );
  MUX2_X1 U4869 ( .A(reg_mem[1272]), .B(reg_mem[1264]), .S(n6770), .Z(n4818)
         );
  MUX2_X1 U4870 ( .A(n4818), .B(n4817), .S(n6719), .Z(n4819) );
  MUX2_X1 U4871 ( .A(n4819), .B(n4816), .S(n6711), .Z(n4820) );
  MUX2_X1 U4872 ( .A(n4820), .B(n4813), .S(n6701), .Z(n4821) );
  MUX2_X1 U4873 ( .A(n4821), .B(n4806), .S(n6700), .Z(n4822) );
  MUX2_X1 U4874 ( .A(reg_mem[1288]), .B(reg_mem[1280]), .S(n6763), .Z(n4823)
         );
  MUX2_X1 U4875 ( .A(reg_mem[1304]), .B(reg_mem[1296]), .S(n6783), .Z(n4824)
         );
  MUX2_X1 U4876 ( .A(n4824), .B(n4823), .S(n6719), .Z(n4825) );
  MUX2_X1 U4877 ( .A(reg_mem[1320]), .B(reg_mem[1312]), .S(n6783), .Z(n4826)
         );
  MUX2_X1 U4878 ( .A(reg_mem[1336]), .B(reg_mem[1328]), .S(n6774), .Z(n4827)
         );
  MUX2_X1 U4879 ( .A(n4827), .B(n4826), .S(n6736), .Z(n4828) );
  MUX2_X1 U4880 ( .A(n4828), .B(n4825), .S(n6716), .Z(n4829) );
  MUX2_X1 U4881 ( .A(reg_mem[1352]), .B(reg_mem[1344]), .S(n6766), .Z(n4830)
         );
  MUX2_X1 U4882 ( .A(reg_mem[1368]), .B(reg_mem[1360]), .S(n6762), .Z(n4831)
         );
  MUX2_X1 U4883 ( .A(n4831), .B(n4830), .S(n6728), .Z(n4832) );
  MUX2_X1 U4884 ( .A(reg_mem[1384]), .B(reg_mem[1376]), .S(n6783), .Z(n4833)
         );
  MUX2_X1 U4885 ( .A(reg_mem[1400]), .B(reg_mem[1392]), .S(n6783), .Z(n4834)
         );
  MUX2_X1 U4886 ( .A(n4834), .B(n4833), .S(n6738), .Z(n4835) );
  MUX2_X1 U4887 ( .A(n4835), .B(n4832), .S(n6715), .Z(n4836) );
  MUX2_X1 U4888 ( .A(n4836), .B(n4829), .S(addr_r[3]), .Z(n4837) );
  MUX2_X1 U4889 ( .A(reg_mem[1416]), .B(reg_mem[1408]), .S(n6748), .Z(n4838)
         );
  MUX2_X1 U4890 ( .A(reg_mem[1432]), .B(reg_mem[1424]), .S(n6772), .Z(n4839)
         );
  MUX2_X1 U4891 ( .A(n4839), .B(n4838), .S(n6732), .Z(n4840) );
  MUX2_X1 U4892 ( .A(reg_mem[1448]), .B(reg_mem[1440]), .S(n6783), .Z(n4841)
         );
  MUX2_X1 U4893 ( .A(reg_mem[1464]), .B(reg_mem[1456]), .S(n6746), .Z(n4842)
         );
  MUX2_X1 U4894 ( .A(n4842), .B(n4841), .S(n6719), .Z(n4843) );
  MUX2_X1 U4895 ( .A(n4843), .B(n4840), .S(n6709), .Z(n4844) );
  MUX2_X1 U4896 ( .A(reg_mem[1480]), .B(reg_mem[1472]), .S(n6775), .Z(n4845)
         );
  MUX2_X1 U4897 ( .A(reg_mem[1496]), .B(reg_mem[1488]), .S(n6777), .Z(n4846)
         );
  MUX2_X1 U4898 ( .A(n4846), .B(n4845), .S(n6725), .Z(n4847) );
  MUX2_X1 U4899 ( .A(reg_mem[1512]), .B(reg_mem[1504]), .S(n6774), .Z(n4848)
         );
  MUX2_X1 U4900 ( .A(reg_mem[1528]), .B(reg_mem[1520]), .S(n6780), .Z(n4849)
         );
  MUX2_X1 U4901 ( .A(n4849), .B(n4848), .S(n6720), .Z(n4850) );
  MUX2_X1 U4902 ( .A(n4850), .B(n4847), .S(addr_r[2]), .Z(n4851) );
  MUX2_X1 U4903 ( .A(n4851), .B(n4844), .S(n6704), .Z(n4852) );
  MUX2_X1 U4904 ( .A(n4852), .B(n4837), .S(n6700), .Z(n4853) );
  MUX2_X1 U4905 ( .A(n4853), .B(n4822), .S(addr_r[5]), .Z(n4854) );
  MUX2_X1 U4906 ( .A(reg_mem[1544]), .B(reg_mem[1536]), .S(n6746), .Z(n4855)
         );
  MUX2_X1 U4907 ( .A(reg_mem[1560]), .B(reg_mem[1552]), .S(n6770), .Z(n4856)
         );
  MUX2_X1 U4908 ( .A(n4856), .B(n4855), .S(n6739), .Z(n4857) );
  MUX2_X1 U4909 ( .A(reg_mem[1576]), .B(reg_mem[1568]), .S(addr_r[0]), .Z(
        n4858) );
  MUX2_X1 U4910 ( .A(reg_mem[1592]), .B(reg_mem[1584]), .S(n6742), .Z(n4859)
         );
  MUX2_X1 U4911 ( .A(n4859), .B(n4858), .S(n6729), .Z(n4860) );
  MUX2_X1 U4912 ( .A(n4860), .B(n4857), .S(n6710), .Z(n4861) );
  MUX2_X1 U4913 ( .A(reg_mem[1608]), .B(reg_mem[1600]), .S(n6761), .Z(n4862)
         );
  MUX2_X1 U4914 ( .A(reg_mem[1624]), .B(reg_mem[1616]), .S(n6763), .Z(n4863)
         );
  MUX2_X1 U4915 ( .A(n4863), .B(n4862), .S(n6724), .Z(n4864) );
  MUX2_X1 U4916 ( .A(reg_mem[1640]), .B(reg_mem[1632]), .S(n6740), .Z(n4865)
         );
  MUX2_X1 U4917 ( .A(reg_mem[1656]), .B(reg_mem[1648]), .S(n6783), .Z(n4866)
         );
  MUX2_X1 U4918 ( .A(n4866), .B(n4865), .S(n6737), .Z(n4867) );
  MUX2_X1 U4919 ( .A(n4867), .B(n4864), .S(n6717), .Z(n4868) );
  MUX2_X1 U4920 ( .A(n4868), .B(n4861), .S(addr_r[3]), .Z(n4869) );
  MUX2_X1 U4921 ( .A(reg_mem[1672]), .B(reg_mem[1664]), .S(n6773), .Z(n4870)
         );
  MUX2_X1 U4922 ( .A(reg_mem[1688]), .B(reg_mem[1680]), .S(n6740), .Z(n4871)
         );
  MUX2_X1 U4923 ( .A(n4871), .B(n4870), .S(n6720), .Z(n4872) );
  MUX2_X1 U4924 ( .A(reg_mem[1704]), .B(reg_mem[1696]), .S(n6783), .Z(n4873)
         );
  MUX2_X1 U4925 ( .A(reg_mem[1720]), .B(reg_mem[1712]), .S(n6759), .Z(n4874)
         );
  MUX2_X1 U4926 ( .A(n4874), .B(n4873), .S(n6731), .Z(n4875) );
  MUX2_X1 U4927 ( .A(n4875), .B(n4872), .S(n6713), .Z(n4876) );
  MUX2_X1 U4928 ( .A(reg_mem[1736]), .B(reg_mem[1728]), .S(n6759), .Z(n4877)
         );
  MUX2_X1 U4929 ( .A(reg_mem[1752]), .B(reg_mem[1744]), .S(n6783), .Z(n4878)
         );
  MUX2_X1 U4930 ( .A(n4878), .B(n4877), .S(n6736), .Z(n4879) );
  MUX2_X1 U4931 ( .A(reg_mem[1768]), .B(reg_mem[1760]), .S(n6780), .Z(n4880)
         );
  MUX2_X1 U4932 ( .A(reg_mem[1784]), .B(reg_mem[1776]), .S(addr_r[0]), .Z(
        n4881) );
  MUX2_X1 U4933 ( .A(n4881), .B(n4880), .S(n6731), .Z(n4882) );
  MUX2_X1 U4934 ( .A(n4882), .B(n4879), .S(addr_r[2]), .Z(n4883) );
  MUX2_X1 U4935 ( .A(n4883), .B(n4876), .S(n6706), .Z(n4884) );
  MUX2_X1 U4936 ( .A(n4884), .B(n4869), .S(n6700), .Z(n4885) );
  MUX2_X1 U4937 ( .A(reg_mem[1800]), .B(reg_mem[1792]), .S(n6746), .Z(n4886)
         );
  MUX2_X1 U4938 ( .A(reg_mem[1816]), .B(reg_mem[1808]), .S(n6776), .Z(n4887)
         );
  MUX2_X1 U4939 ( .A(n4887), .B(n4886), .S(n6723), .Z(n4888) );
  MUX2_X1 U4940 ( .A(reg_mem[1832]), .B(reg_mem[1824]), .S(n6769), .Z(n4889)
         );
  MUX2_X1 U4941 ( .A(reg_mem[1848]), .B(reg_mem[1840]), .S(n6743), .Z(n4890)
         );
  MUX2_X1 U4942 ( .A(n4890), .B(n4889), .S(n6720), .Z(n4891) );
  MUX2_X1 U4943 ( .A(n4891), .B(n4888), .S(n6714), .Z(n4892) );
  MUX2_X1 U4944 ( .A(reg_mem[1864]), .B(reg_mem[1856]), .S(n6747), .Z(n4893)
         );
  MUX2_X1 U4945 ( .A(reg_mem[1880]), .B(reg_mem[1872]), .S(n6745), .Z(n4894)
         );
  MUX2_X1 U4946 ( .A(n4894), .B(n4893), .S(n6736), .Z(n4895) );
  MUX2_X1 U4947 ( .A(reg_mem[1896]), .B(reg_mem[1888]), .S(n6774), .Z(n4896)
         );
  MUX2_X1 U4948 ( .A(reg_mem[1912]), .B(reg_mem[1904]), .S(n6779), .Z(n4897)
         );
  MUX2_X1 U4949 ( .A(n4897), .B(n4896), .S(n6719), .Z(n4898) );
  MUX2_X1 U4950 ( .A(n4898), .B(n4895), .S(n6708), .Z(n4899) );
  MUX2_X1 U4951 ( .A(n4899), .B(n4892), .S(n6706), .Z(n4900) );
  MUX2_X1 U4952 ( .A(reg_mem[1928]), .B(reg_mem[1920]), .S(n6764), .Z(n4901)
         );
  MUX2_X1 U4953 ( .A(reg_mem[1944]), .B(reg_mem[1936]), .S(n6750), .Z(n4902)
         );
  MUX2_X1 U4954 ( .A(n4902), .B(n4901), .S(n6726), .Z(n4903) );
  MUX2_X1 U4955 ( .A(reg_mem[1960]), .B(reg_mem[1952]), .S(n6756), .Z(n4904)
         );
  MUX2_X1 U4956 ( .A(reg_mem[1976]), .B(reg_mem[1968]), .S(n6775), .Z(n4905)
         );
  MUX2_X1 U4957 ( .A(n4905), .B(n4904), .S(n6719), .Z(n4906) );
  MUX2_X1 U4958 ( .A(n4906), .B(n4903), .S(n6708), .Z(n4907) );
  MUX2_X1 U4959 ( .A(reg_mem[1992]), .B(reg_mem[1984]), .S(n6741), .Z(n4908)
         );
  MUX2_X1 U4960 ( .A(reg_mem[2008]), .B(reg_mem[2000]), .S(n6740), .Z(n4909)
         );
  MUX2_X1 U4961 ( .A(n4909), .B(n4908), .S(n6737), .Z(n4910) );
  MUX2_X1 U4962 ( .A(reg_mem[2024]), .B(reg_mem[2016]), .S(n6769), .Z(n4911)
         );
  MUX2_X1 U4963 ( .A(reg_mem[2040]), .B(reg_mem[2032]), .S(n6741), .Z(n4912)
         );
  MUX2_X1 U4964 ( .A(n4912), .B(n4911), .S(n6731), .Z(n4913) );
  MUX2_X1 U4965 ( .A(n4913), .B(n4910), .S(n6710), .Z(n4914) );
  MUX2_X1 U4966 ( .A(n4914), .B(n4907), .S(n6703), .Z(n4915) );
  MUX2_X1 U4967 ( .A(n4915), .B(n4900), .S(n6700), .Z(n4916) );
  MUX2_X1 U4968 ( .A(n4916), .B(n4885), .S(addr_r[5]), .Z(n4917) );
  MUX2_X1 U4969 ( .A(n4917), .B(n4854), .S(addr_r[6]), .Z(n4918) );
  MUX2_X1 U4970 ( .A(n4918), .B(n4791), .S(addr_r[7]), .Z(data_r[0]) );
  MUX2_X1 U4971 ( .A(reg_mem[9]), .B(reg_mem[1]), .S(n6742), .Z(n4919) );
  MUX2_X1 U4972 ( .A(reg_mem[25]), .B(reg_mem[17]), .S(n6777), .Z(n4920) );
  MUX2_X1 U4973 ( .A(n4920), .B(n4919), .S(n6720), .Z(n4921) );
  MUX2_X1 U4974 ( .A(reg_mem[41]), .B(reg_mem[33]), .S(n6764), .Z(n4922) );
  MUX2_X1 U4975 ( .A(reg_mem[57]), .B(reg_mem[49]), .S(n6749), .Z(n4923) );
  MUX2_X1 U4976 ( .A(n4923), .B(n4922), .S(n6724), .Z(n4924) );
  MUX2_X1 U4977 ( .A(n4924), .B(n4921), .S(n6708), .Z(n4925) );
  MUX2_X1 U4978 ( .A(reg_mem[73]), .B(reg_mem[65]), .S(n6759), .Z(n4926) );
  MUX2_X1 U4979 ( .A(reg_mem[89]), .B(reg_mem[81]), .S(n6758), .Z(n4927) );
  MUX2_X1 U4980 ( .A(n4927), .B(n4926), .S(n6719), .Z(n4928) );
  MUX2_X1 U4981 ( .A(reg_mem[105]), .B(reg_mem[97]), .S(n6745), .Z(n4929) );
  MUX2_X1 U4982 ( .A(reg_mem[121]), .B(reg_mem[113]), .S(n6741), .Z(n4930) );
  MUX2_X1 U4983 ( .A(n4930), .B(n4929), .S(n6719), .Z(n4931) );
  MUX2_X1 U4984 ( .A(n4931), .B(n4928), .S(n6717), .Z(n4932) );
  MUX2_X1 U4985 ( .A(n4932), .B(n4925), .S(n6701), .Z(n4933) );
  MUX2_X1 U4986 ( .A(reg_mem[137]), .B(reg_mem[129]), .S(n6778), .Z(n4934) );
  MUX2_X1 U4987 ( .A(reg_mem[153]), .B(reg_mem[145]), .S(n6740), .Z(n4935) );
  MUX2_X1 U4988 ( .A(n4935), .B(n4934), .S(n6718), .Z(n4936) );
  MUX2_X1 U4989 ( .A(reg_mem[169]), .B(reg_mem[161]), .S(n6748), .Z(n4937) );
  MUX2_X1 U4990 ( .A(reg_mem[185]), .B(reg_mem[177]), .S(n6758), .Z(n4938) );
  MUX2_X1 U4991 ( .A(n4938), .B(n4937), .S(n6718), .Z(n4939) );
  MUX2_X1 U4992 ( .A(n4939), .B(n4936), .S(n6712), .Z(n4940) );
  MUX2_X1 U4993 ( .A(reg_mem[201]), .B(reg_mem[193]), .S(n6741), .Z(n4941) );
  MUX2_X1 U4994 ( .A(reg_mem[217]), .B(reg_mem[209]), .S(n6742), .Z(n4942) );
  MUX2_X1 U4995 ( .A(n4942), .B(n4941), .S(n6723), .Z(n4943) );
  MUX2_X1 U4996 ( .A(reg_mem[233]), .B(reg_mem[225]), .S(n6783), .Z(n4944) );
  MUX2_X1 U4997 ( .A(reg_mem[249]), .B(reg_mem[241]), .S(n6783), .Z(n4945) );
  MUX2_X1 U4998 ( .A(n4945), .B(n4944), .S(n6739), .Z(n4946) );
  MUX2_X1 U4999 ( .A(n4946), .B(n4943), .S(n6717), .Z(n4947) );
  MUX2_X1 U5000 ( .A(n4947), .B(n4940), .S(n6704), .Z(n4948) );
  MUX2_X1 U5001 ( .A(n4948), .B(n4933), .S(n6700), .Z(n4949) );
  MUX2_X1 U5002 ( .A(reg_mem[265]), .B(reg_mem[257]), .S(n6779), .Z(n4950) );
  MUX2_X1 U5003 ( .A(reg_mem[281]), .B(reg_mem[273]), .S(n6758), .Z(n4951) );
  MUX2_X1 U5004 ( .A(n4951), .B(n4950), .S(n6718), .Z(n4952) );
  MUX2_X1 U5005 ( .A(reg_mem[297]), .B(reg_mem[289]), .S(n6742), .Z(n4953) );
  MUX2_X1 U5006 ( .A(reg_mem[313]), .B(reg_mem[305]), .S(n6753), .Z(n4954) );
  MUX2_X1 U5007 ( .A(n4954), .B(n4953), .S(n6724), .Z(n4955) );
  MUX2_X1 U5008 ( .A(n4955), .B(n4952), .S(n6716), .Z(n4956) );
  MUX2_X1 U5009 ( .A(reg_mem[329]), .B(reg_mem[321]), .S(n6742), .Z(n4957) );
  MUX2_X1 U5010 ( .A(reg_mem[345]), .B(reg_mem[337]), .S(n6770), .Z(n4958) );
  MUX2_X1 U5011 ( .A(n4958), .B(n4957), .S(n6722), .Z(n4959) );
  MUX2_X1 U5012 ( .A(reg_mem[361]), .B(reg_mem[353]), .S(n6759), .Z(n4960) );
  MUX2_X1 U5013 ( .A(reg_mem[377]), .B(reg_mem[369]), .S(n6767), .Z(n4961) );
  MUX2_X1 U5014 ( .A(n4961), .B(n4960), .S(n6724), .Z(n4962) );
  MUX2_X1 U5015 ( .A(n4962), .B(n4959), .S(n6713), .Z(n4963) );
  MUX2_X1 U5016 ( .A(n4963), .B(n4956), .S(n6703), .Z(n4964) );
  MUX2_X1 U5017 ( .A(reg_mem[393]), .B(reg_mem[385]), .S(n6764), .Z(n4965) );
  MUX2_X1 U5018 ( .A(reg_mem[409]), .B(reg_mem[401]), .S(n6741), .Z(n4966) );
  MUX2_X1 U5019 ( .A(n4966), .B(n4965), .S(n6718), .Z(n4967) );
  MUX2_X1 U5020 ( .A(reg_mem[425]), .B(reg_mem[417]), .S(n6756), .Z(n4968) );
  MUX2_X1 U5021 ( .A(reg_mem[441]), .B(reg_mem[433]), .S(n6759), .Z(n4969) );
  MUX2_X1 U5022 ( .A(n4969), .B(n4968), .S(n6721), .Z(n4970) );
  MUX2_X1 U5023 ( .A(n4970), .B(n4967), .S(addr_r[2]), .Z(n4971) );
  MUX2_X1 U5024 ( .A(reg_mem[457]), .B(reg_mem[449]), .S(n6778), .Z(n4972) );
  MUX2_X1 U5025 ( .A(reg_mem[473]), .B(reg_mem[465]), .S(n6742), .Z(n4973) );
  MUX2_X1 U5026 ( .A(n4973), .B(n4972), .S(n6718), .Z(n4974) );
  MUX2_X1 U5027 ( .A(reg_mem[489]), .B(reg_mem[481]), .S(n6760), .Z(n4975) );
  MUX2_X1 U5028 ( .A(reg_mem[505]), .B(reg_mem[497]), .S(n6759), .Z(n4976) );
  MUX2_X1 U5029 ( .A(n4976), .B(n4975), .S(n6720), .Z(n4977) );
  MUX2_X1 U5030 ( .A(n4977), .B(n4974), .S(n6708), .Z(n4978) );
  MUX2_X1 U5031 ( .A(n4978), .B(n4971), .S(n6702), .Z(n4979) );
  MUX2_X1 U5032 ( .A(n4979), .B(n4964), .S(n6700), .Z(n4980) );
  MUX2_X1 U5033 ( .A(n4980), .B(n4949), .S(n6697), .Z(n4981) );
  MUX2_X1 U5034 ( .A(reg_mem[521]), .B(reg_mem[513]), .S(n6758), .Z(n4982) );
  MUX2_X1 U5035 ( .A(reg_mem[537]), .B(reg_mem[529]), .S(n6756), .Z(n4983) );
  MUX2_X1 U5036 ( .A(n4983), .B(n4982), .S(n6720), .Z(n4984) );
  MUX2_X1 U5037 ( .A(reg_mem[553]), .B(reg_mem[545]), .S(n6741), .Z(n4985) );
  MUX2_X1 U5038 ( .A(reg_mem[569]), .B(reg_mem[561]), .S(n6740), .Z(n4986) );
  MUX2_X1 U5039 ( .A(n4986), .B(n4985), .S(n6739), .Z(n4987) );
  MUX2_X1 U5040 ( .A(n4987), .B(n4984), .S(n6714), .Z(n4988) );
  MUX2_X1 U5041 ( .A(reg_mem[585]), .B(reg_mem[577]), .S(n6742), .Z(n4989) );
  MUX2_X1 U5042 ( .A(reg_mem[601]), .B(reg_mem[593]), .S(n6742), .Z(n4990) );
  MUX2_X1 U5043 ( .A(n4990), .B(n4989), .S(n6720), .Z(n4991) );
  MUX2_X1 U5044 ( .A(reg_mem[617]), .B(reg_mem[609]), .S(n6767), .Z(n4992) );
  MUX2_X1 U5045 ( .A(reg_mem[633]), .B(reg_mem[625]), .S(n6740), .Z(n4993) );
  MUX2_X1 U5046 ( .A(n4993), .B(n4992), .S(n6739), .Z(n4994) );
  MUX2_X1 U5047 ( .A(n4994), .B(n4991), .S(n6709), .Z(n4995) );
  MUX2_X1 U5048 ( .A(n4995), .B(n4988), .S(n6705), .Z(n4996) );
  MUX2_X1 U5049 ( .A(reg_mem[649]), .B(reg_mem[641]), .S(n6740), .Z(n4997) );
  MUX2_X1 U5050 ( .A(reg_mem[665]), .B(reg_mem[657]), .S(n6761), .Z(n4998) );
  MUX2_X1 U5051 ( .A(n4998), .B(n4997), .S(n6726), .Z(n4999) );
  MUX2_X1 U5052 ( .A(reg_mem[681]), .B(reg_mem[673]), .S(n6754), .Z(n5000) );
  MUX2_X1 U5053 ( .A(reg_mem[697]), .B(reg_mem[689]), .S(n6741), .Z(n5001) );
  MUX2_X1 U5054 ( .A(n5001), .B(n5000), .S(n6738), .Z(n5002) );
  MUX2_X1 U5055 ( .A(n5002), .B(n4999), .S(n6714), .Z(n5003) );
  MUX2_X1 U5056 ( .A(reg_mem[713]), .B(reg_mem[705]), .S(n6743), .Z(n5004) );
  MUX2_X1 U5057 ( .A(reg_mem[729]), .B(reg_mem[721]), .S(n6751), .Z(n5005) );
  MUX2_X1 U5058 ( .A(n5005), .B(n5004), .S(n6718), .Z(n5006) );
  MUX2_X1 U5059 ( .A(reg_mem[745]), .B(reg_mem[737]), .S(n6761), .Z(n5007) );
  MUX2_X1 U5060 ( .A(reg_mem[761]), .B(reg_mem[753]), .S(n6781), .Z(n5008) );
  MUX2_X1 U5061 ( .A(n5008), .B(n5007), .S(n6739), .Z(n5009) );
  MUX2_X1 U5062 ( .A(n5009), .B(n5006), .S(n6707), .Z(n5010) );
  MUX2_X1 U5063 ( .A(n5010), .B(n5003), .S(n6706), .Z(n5011) );
  MUX2_X1 U5064 ( .A(n5011), .B(n4996), .S(n6700), .Z(n5012) );
  MUX2_X1 U5065 ( .A(reg_mem[777]), .B(reg_mem[769]), .S(n6747), .Z(n5013) );
  MUX2_X1 U5066 ( .A(reg_mem[793]), .B(reg_mem[785]), .S(n6774), .Z(n5014) );
  MUX2_X1 U5067 ( .A(n5014), .B(n5013), .S(n6718), .Z(n5015) );
  MUX2_X1 U5068 ( .A(reg_mem[809]), .B(reg_mem[801]), .S(n6780), .Z(n5016) );
  MUX2_X1 U5069 ( .A(reg_mem[825]), .B(reg_mem[817]), .S(n6747), .Z(n5017) );
  MUX2_X1 U5070 ( .A(n5017), .B(n5016), .S(n6721), .Z(n5018) );
  MUX2_X1 U5071 ( .A(n5018), .B(n5015), .S(n6716), .Z(n5019) );
  MUX2_X1 U5072 ( .A(reg_mem[841]), .B(reg_mem[833]), .S(n6776), .Z(n5020) );
  MUX2_X1 U5073 ( .A(reg_mem[857]), .B(reg_mem[849]), .S(n6750), .Z(n5021) );
  MUX2_X1 U5074 ( .A(n5021), .B(n5020), .S(n6721), .Z(n5022) );
  MUX2_X1 U5075 ( .A(reg_mem[873]), .B(reg_mem[865]), .S(n6748), .Z(n5023) );
  MUX2_X1 U5076 ( .A(reg_mem[889]), .B(reg_mem[881]), .S(n6767), .Z(n5024) );
  MUX2_X1 U5077 ( .A(n5024), .B(n5023), .S(n6727), .Z(n5025) );
  MUX2_X1 U5078 ( .A(n5025), .B(n5022), .S(n6715), .Z(n5026) );
  MUX2_X1 U5079 ( .A(n5026), .B(n5019), .S(n6702), .Z(n5027) );
  MUX2_X1 U5080 ( .A(reg_mem[905]), .B(reg_mem[897]), .S(n6754), .Z(n5028) );
  MUX2_X1 U5081 ( .A(reg_mem[921]), .B(reg_mem[913]), .S(n6757), .Z(n5029) );
  MUX2_X1 U5082 ( .A(n5029), .B(n5028), .S(n6724), .Z(n5030) );
  MUX2_X1 U5083 ( .A(reg_mem[937]), .B(reg_mem[929]), .S(n6758), .Z(n5031) );
  MUX2_X1 U5084 ( .A(reg_mem[953]), .B(reg_mem[945]), .S(n6762), .Z(n5032) );
  MUX2_X1 U5085 ( .A(n5032), .B(n5031), .S(n6735), .Z(n5033) );
  MUX2_X1 U5086 ( .A(n5033), .B(n5030), .S(n6710), .Z(n5034) );
  MUX2_X1 U5087 ( .A(reg_mem[969]), .B(reg_mem[961]), .S(n6750), .Z(n5035) );
  MUX2_X1 U5088 ( .A(reg_mem[985]), .B(reg_mem[977]), .S(n6767), .Z(n5036) );
  MUX2_X1 U5089 ( .A(n5036), .B(n5035), .S(n6721), .Z(n5037) );
  MUX2_X1 U5090 ( .A(reg_mem[1001]), .B(reg_mem[993]), .S(n6752), .Z(n5038) );
  MUX2_X1 U5091 ( .A(reg_mem[1017]), .B(reg_mem[1009]), .S(n6768), .Z(n5039)
         );
  MUX2_X1 U5092 ( .A(n5039), .B(n5038), .S(n6734), .Z(n5040) );
  MUX2_X1 U5093 ( .A(n5040), .B(n5037), .S(n6714), .Z(n5041) );
  MUX2_X1 U5094 ( .A(n5041), .B(n5034), .S(n6704), .Z(n5042) );
  MUX2_X1 U5095 ( .A(n5042), .B(n5027), .S(n6700), .Z(n5043) );
  MUX2_X1 U5096 ( .A(n5043), .B(n5012), .S(addr_r[5]), .Z(n5044) );
  MUX2_X1 U5097 ( .A(n5044), .B(n4981), .S(addr_r[6]), .Z(n5045) );
  MUX2_X1 U5098 ( .A(reg_mem[1033]), .B(reg_mem[1025]), .S(n6765), .Z(n5046)
         );
  MUX2_X1 U5099 ( .A(reg_mem[1049]), .B(reg_mem[1041]), .S(n6749), .Z(n5047)
         );
  MUX2_X1 U5100 ( .A(n5047), .B(n5046), .S(n6733), .Z(n5048) );
  MUX2_X1 U5101 ( .A(reg_mem[1065]), .B(reg_mem[1057]), .S(n6748), .Z(n5049)
         );
  MUX2_X1 U5102 ( .A(reg_mem[1081]), .B(reg_mem[1073]), .S(n6780), .Z(n5050)
         );
  MUX2_X1 U5103 ( .A(n5050), .B(n5049), .S(n6739), .Z(n5051) );
  MUX2_X1 U5104 ( .A(n5051), .B(n5048), .S(n6709), .Z(n5052) );
  MUX2_X1 U5105 ( .A(reg_mem[1097]), .B(reg_mem[1089]), .S(n6772), .Z(n5053)
         );
  MUX2_X1 U5106 ( .A(reg_mem[1113]), .B(reg_mem[1105]), .S(n6774), .Z(n5054)
         );
  MUX2_X1 U5107 ( .A(n5054), .B(n5053), .S(n6725), .Z(n5055) );
  MUX2_X1 U5108 ( .A(reg_mem[1129]), .B(reg_mem[1121]), .S(n6773), .Z(n5056)
         );
  MUX2_X1 U5109 ( .A(reg_mem[1145]), .B(reg_mem[1137]), .S(n6768), .Z(n5057)
         );
  MUX2_X1 U5110 ( .A(n5057), .B(n5056), .S(n6737), .Z(n5058) );
  MUX2_X1 U5111 ( .A(n5058), .B(n5055), .S(n6716), .Z(n5059) );
  MUX2_X1 U5112 ( .A(n5059), .B(n5052), .S(n6705), .Z(n5060) );
  MUX2_X1 U5113 ( .A(reg_mem[1161]), .B(reg_mem[1153]), .S(n6765), .Z(n5061)
         );
  MUX2_X1 U5114 ( .A(reg_mem[1177]), .B(reg_mem[1169]), .S(n6776), .Z(n5062)
         );
  MUX2_X1 U5115 ( .A(n5062), .B(n5061), .S(n6728), .Z(n5063) );
  MUX2_X1 U5116 ( .A(reg_mem[1193]), .B(reg_mem[1185]), .S(n6766), .Z(n5064)
         );
  MUX2_X1 U5117 ( .A(reg_mem[1209]), .B(reg_mem[1201]), .S(n6767), .Z(n5065)
         );
  MUX2_X1 U5118 ( .A(n5065), .B(n5064), .S(n6732), .Z(n5066) );
  MUX2_X1 U5119 ( .A(n5066), .B(n5063), .S(n6712), .Z(n5067) );
  MUX2_X1 U5120 ( .A(reg_mem[1225]), .B(reg_mem[1217]), .S(n6763), .Z(n5068)
         );
  MUX2_X1 U5121 ( .A(reg_mem[1241]), .B(reg_mem[1233]), .S(n6769), .Z(n5069)
         );
  MUX2_X1 U5122 ( .A(n5069), .B(n5068), .S(n6722), .Z(n5070) );
  MUX2_X1 U5123 ( .A(reg_mem[1257]), .B(reg_mem[1249]), .S(n6771), .Z(n5071)
         );
  MUX2_X1 U5124 ( .A(reg_mem[1273]), .B(reg_mem[1265]), .S(n6761), .Z(n5072)
         );
  MUX2_X1 U5125 ( .A(n5072), .B(n5071), .S(n6737), .Z(n5073) );
  MUX2_X1 U5126 ( .A(n5073), .B(n5070), .S(n6711), .Z(n5074) );
  MUX2_X1 U5127 ( .A(n5074), .B(n5067), .S(n6706), .Z(n5075) );
  MUX2_X1 U5128 ( .A(n5075), .B(n5060), .S(n6700), .Z(n5076) );
  MUX2_X1 U5129 ( .A(reg_mem[1289]), .B(reg_mem[1281]), .S(n6777), .Z(n5077)
         );
  MUX2_X1 U5130 ( .A(reg_mem[1305]), .B(reg_mem[1297]), .S(n6755), .Z(n5078)
         );
  MUX2_X1 U5131 ( .A(n5078), .B(n5077), .S(n6721), .Z(n5079) );
  MUX2_X1 U5132 ( .A(reg_mem[1321]), .B(reg_mem[1313]), .S(n6771), .Z(n5080)
         );
  MUX2_X1 U5133 ( .A(reg_mem[1337]), .B(reg_mem[1329]), .S(n6741), .Z(n5081)
         );
  MUX2_X1 U5134 ( .A(n5081), .B(n5080), .S(n6720), .Z(n5082) );
  MUX2_X1 U5135 ( .A(n5082), .B(n5079), .S(n6707), .Z(n5083) );
  MUX2_X1 U5136 ( .A(reg_mem[1353]), .B(reg_mem[1345]), .S(n6773), .Z(n5084)
         );
  MUX2_X1 U5137 ( .A(reg_mem[1369]), .B(reg_mem[1361]), .S(n6759), .Z(n5085)
         );
  MUX2_X1 U5138 ( .A(n5085), .B(n5084), .S(n6728), .Z(n5086) );
  MUX2_X1 U5139 ( .A(reg_mem[1385]), .B(reg_mem[1377]), .S(n6751), .Z(n5087)
         );
  MUX2_X1 U5140 ( .A(reg_mem[1401]), .B(reg_mem[1393]), .S(n6783), .Z(n5088)
         );
  MUX2_X1 U5141 ( .A(n5088), .B(n5087), .S(n6727), .Z(n5089) );
  MUX2_X1 U5142 ( .A(n5089), .B(n5086), .S(n6713), .Z(n5090) );
  MUX2_X1 U5143 ( .A(n5090), .B(n5083), .S(n6703), .Z(n5091) );
  MUX2_X1 U5144 ( .A(reg_mem[1417]), .B(reg_mem[1409]), .S(n6758), .Z(n5092)
         );
  MUX2_X1 U5145 ( .A(reg_mem[1433]), .B(reg_mem[1425]), .S(n6742), .Z(n5093)
         );
  MUX2_X1 U5146 ( .A(n5093), .B(n5092), .S(n6726), .Z(n5094) );
  MUX2_X1 U5147 ( .A(reg_mem[1449]), .B(reg_mem[1441]), .S(n6740), .Z(n5095)
         );
  MUX2_X1 U5148 ( .A(reg_mem[1465]), .B(reg_mem[1457]), .S(n6740), .Z(n5096)
         );
  MUX2_X1 U5149 ( .A(n5096), .B(n5095), .S(n6732), .Z(n5097) );
  MUX2_X1 U5150 ( .A(n5097), .B(n5094), .S(n6710), .Z(n5098) );
  MUX2_X1 U5151 ( .A(reg_mem[1481]), .B(reg_mem[1473]), .S(n6761), .Z(n5099)
         );
  MUX2_X1 U5152 ( .A(reg_mem[1497]), .B(reg_mem[1489]), .S(n6766), .Z(n5100)
         );
  MUX2_X1 U5153 ( .A(n5100), .B(n5099), .S(n6731), .Z(n5101) );
  MUX2_X1 U5154 ( .A(reg_mem[1513]), .B(reg_mem[1505]), .S(n6778), .Z(n5102)
         );
  MUX2_X1 U5155 ( .A(reg_mem[1529]), .B(reg_mem[1521]), .S(n6740), .Z(n5103)
         );
  MUX2_X1 U5156 ( .A(n5103), .B(n5102), .S(n6719), .Z(n5104) );
  MUX2_X1 U5157 ( .A(n5104), .B(n5101), .S(n6714), .Z(n5105) );
  MUX2_X1 U5158 ( .A(n5105), .B(n5098), .S(n6701), .Z(n5106) );
  MUX2_X1 U5159 ( .A(n5106), .B(n5091), .S(n6700), .Z(n5107) );
  MUX2_X1 U5160 ( .A(n5107), .B(n5076), .S(addr_r[5]), .Z(n5108) );
  MUX2_X1 U5161 ( .A(reg_mem[1545]), .B(reg_mem[1537]), .S(n6776), .Z(n5109)
         );
  MUX2_X1 U5162 ( .A(reg_mem[1561]), .B(reg_mem[1553]), .S(n6742), .Z(n5110)
         );
  MUX2_X1 U5163 ( .A(n5110), .B(n5109), .S(n6732), .Z(n5111) );
  MUX2_X1 U5164 ( .A(reg_mem[1577]), .B(reg_mem[1569]), .S(n6740), .Z(n5112)
         );
  MUX2_X1 U5165 ( .A(reg_mem[1593]), .B(reg_mem[1585]), .S(n6773), .Z(n5113)
         );
  MUX2_X1 U5166 ( .A(n5113), .B(n5112), .S(n6726), .Z(n5114) );
  MUX2_X1 U5167 ( .A(n5114), .B(n5111), .S(n6707), .Z(n5115) );
  MUX2_X1 U5168 ( .A(reg_mem[1609]), .B(reg_mem[1601]), .S(n6783), .Z(n5116)
         );
  MUX2_X1 U5169 ( .A(reg_mem[1625]), .B(reg_mem[1617]), .S(n6750), .Z(n5117)
         );
  MUX2_X1 U5170 ( .A(n5117), .B(n5116), .S(n6718), .Z(n5118) );
  MUX2_X1 U5171 ( .A(reg_mem[1641]), .B(reg_mem[1633]), .S(n6782), .Z(n5119)
         );
  MUX2_X1 U5172 ( .A(reg_mem[1657]), .B(reg_mem[1649]), .S(addr_r[0]), .Z(
        n5120) );
  MUX2_X1 U5173 ( .A(n5120), .B(n5119), .S(n6733), .Z(n5121) );
  MUX2_X1 U5174 ( .A(n5121), .B(n5118), .S(n6708), .Z(n5122) );
  MUX2_X1 U5175 ( .A(n5122), .B(n5115), .S(n6701), .Z(n5123) );
  MUX2_X1 U5176 ( .A(reg_mem[1673]), .B(reg_mem[1665]), .S(n6763), .Z(n5124)
         );
  MUX2_X1 U5177 ( .A(reg_mem[1689]), .B(reg_mem[1681]), .S(n6761), .Z(n5125)
         );
  MUX2_X1 U5178 ( .A(n5125), .B(n5124), .S(addr_r[1]), .Z(n5126) );
  MUX2_X1 U5179 ( .A(reg_mem[1705]), .B(reg_mem[1697]), .S(n6758), .Z(n5127)
         );
  MUX2_X1 U5180 ( .A(reg_mem[1721]), .B(reg_mem[1713]), .S(n6771), .Z(n5128)
         );
  MUX2_X1 U5181 ( .A(n5128), .B(n5127), .S(addr_r[1]), .Z(n5129) );
  MUX2_X1 U5182 ( .A(n5129), .B(n5126), .S(n6709), .Z(n5130) );
  MUX2_X1 U5183 ( .A(reg_mem[1737]), .B(reg_mem[1729]), .S(n6742), .Z(n5131)
         );
  MUX2_X1 U5184 ( .A(reg_mem[1753]), .B(reg_mem[1745]), .S(n6771), .Z(n5132)
         );
  MUX2_X1 U5185 ( .A(n5132), .B(n5131), .S(addr_r[1]), .Z(n5133) );
  MUX2_X1 U5186 ( .A(reg_mem[1769]), .B(reg_mem[1761]), .S(n6780), .Z(n5134)
         );
  MUX2_X1 U5187 ( .A(reg_mem[1785]), .B(reg_mem[1777]), .S(n6783), .Z(n5135)
         );
  MUX2_X1 U5188 ( .A(n5135), .B(n5134), .S(n6739), .Z(n5136) );
  MUX2_X1 U5189 ( .A(n5136), .B(n5133), .S(n6708), .Z(n5137) );
  MUX2_X1 U5190 ( .A(n5137), .B(n5130), .S(n6705), .Z(n5138) );
  MUX2_X1 U5191 ( .A(n5138), .B(n5123), .S(n6700), .Z(n5139) );
  MUX2_X1 U5192 ( .A(reg_mem[1801]), .B(reg_mem[1793]), .S(n6769), .Z(n5140)
         );
  MUX2_X1 U5193 ( .A(reg_mem[1817]), .B(reg_mem[1809]), .S(n6780), .Z(n5141)
         );
  MUX2_X1 U5194 ( .A(n5141), .B(n5140), .S(addr_r[1]), .Z(n5142) );
  MUX2_X1 U5195 ( .A(reg_mem[1833]), .B(reg_mem[1825]), .S(n6741), .Z(n5143)
         );
  MUX2_X1 U5196 ( .A(reg_mem[1849]), .B(reg_mem[1841]), .S(n6776), .Z(n5144)
         );
  MUX2_X1 U5197 ( .A(n5144), .B(n5143), .S(addr_r[1]), .Z(n5145) );
  MUX2_X1 U5198 ( .A(n5145), .B(n5142), .S(n6713), .Z(n5146) );
  MUX2_X1 U5199 ( .A(reg_mem[1865]), .B(reg_mem[1857]), .S(n6763), .Z(n5147)
         );
  MUX2_X1 U5200 ( .A(reg_mem[1881]), .B(reg_mem[1873]), .S(n6769), .Z(n5148)
         );
  MUX2_X1 U5201 ( .A(n5148), .B(n5147), .S(n6730), .Z(n5149) );
  MUX2_X1 U5202 ( .A(reg_mem[1897]), .B(reg_mem[1889]), .S(n6765), .Z(n5150)
         );
  MUX2_X1 U5203 ( .A(reg_mem[1913]), .B(reg_mem[1905]), .S(n6776), .Z(n5151)
         );
  MUX2_X1 U5204 ( .A(n5151), .B(n5150), .S(n6736), .Z(n5152) );
  MUX2_X1 U5205 ( .A(n5152), .B(n5149), .S(n6710), .Z(n5153) );
  MUX2_X1 U5206 ( .A(n5153), .B(n5146), .S(n6703), .Z(n5154) );
  MUX2_X1 U5207 ( .A(reg_mem[1929]), .B(reg_mem[1921]), .S(n6770), .Z(n5155)
         );
  MUX2_X1 U5208 ( .A(reg_mem[1945]), .B(reg_mem[1937]), .S(n6742), .Z(n5156)
         );
  MUX2_X1 U5209 ( .A(n5156), .B(n5155), .S(n6726), .Z(n5157) );
  MUX2_X1 U5210 ( .A(reg_mem[1961]), .B(reg_mem[1953]), .S(n6765), .Z(n5158)
         );
  MUX2_X1 U5211 ( .A(reg_mem[1977]), .B(reg_mem[1969]), .S(n6758), .Z(n5159)
         );
  MUX2_X1 U5212 ( .A(n5159), .B(n5158), .S(n6738), .Z(n5160) );
  MUX2_X1 U5213 ( .A(n5160), .B(n5157), .S(n6710), .Z(n5161) );
  MUX2_X1 U5214 ( .A(reg_mem[1993]), .B(reg_mem[1985]), .S(n6783), .Z(n5162)
         );
  MUX2_X1 U5215 ( .A(reg_mem[2009]), .B(reg_mem[2001]), .S(n6741), .Z(n5163)
         );
  MUX2_X1 U5216 ( .A(n5163), .B(n5162), .S(n6739), .Z(n5164) );
  MUX2_X1 U5217 ( .A(reg_mem[2025]), .B(reg_mem[2017]), .S(n6768), .Z(n5165)
         );
  MUX2_X1 U5218 ( .A(reg_mem[2041]), .B(reg_mem[2033]), .S(n6783), .Z(n5166)
         );
  MUX2_X1 U5219 ( .A(n5166), .B(n5165), .S(n6739), .Z(n5167) );
  MUX2_X1 U5220 ( .A(n5167), .B(n5164), .S(n6715), .Z(n5168) );
  MUX2_X1 U5221 ( .A(n5168), .B(n5161), .S(n6702), .Z(n5169) );
  MUX2_X1 U5222 ( .A(n5169), .B(n5154), .S(n6700), .Z(n5170) );
  MUX2_X1 U5223 ( .A(n5170), .B(n5139), .S(addr_r[5]), .Z(n5171) );
  MUX2_X1 U5224 ( .A(n5171), .B(n5108), .S(addr_r[6]), .Z(n5172) );
  MUX2_X1 U5225 ( .A(n5172), .B(n5045), .S(addr_r[7]), .Z(data_r[1]) );
  MUX2_X1 U5226 ( .A(reg_mem[10]), .B(reg_mem[2]), .S(n6773), .Z(n5173) );
  MUX2_X1 U5227 ( .A(reg_mem[26]), .B(reg_mem[18]), .S(n6771), .Z(n5174) );
  MUX2_X1 U5228 ( .A(n5174), .B(n5173), .S(n6718), .Z(n5175) );
  MUX2_X1 U5229 ( .A(reg_mem[42]), .B(reg_mem[34]), .S(n6767), .Z(n5176) );
  MUX2_X1 U5230 ( .A(reg_mem[58]), .B(reg_mem[50]), .S(n6744), .Z(n5177) );
  MUX2_X1 U5231 ( .A(n5177), .B(n5176), .S(n6726), .Z(n5178) );
  MUX2_X1 U5232 ( .A(n5178), .B(n5175), .S(n6717), .Z(n5179) );
  MUX2_X1 U5233 ( .A(reg_mem[74]), .B(reg_mem[66]), .S(n6769), .Z(n5180) );
  MUX2_X1 U5234 ( .A(reg_mem[90]), .B(reg_mem[82]), .S(n6778), .Z(n5181) );
  MUX2_X1 U5235 ( .A(n5181), .B(n5180), .S(n6722), .Z(n5182) );
  MUX2_X1 U5236 ( .A(reg_mem[106]), .B(reg_mem[98]), .S(n6782), .Z(n5183) );
  MUX2_X1 U5237 ( .A(reg_mem[122]), .B(reg_mem[114]), .S(n6777), .Z(n5184) );
  MUX2_X1 U5238 ( .A(n5184), .B(n5183), .S(n6721), .Z(n5185) );
  MUX2_X1 U5239 ( .A(n5185), .B(n5182), .S(n6717), .Z(n5186) );
  MUX2_X1 U5240 ( .A(n5186), .B(n5179), .S(n6701), .Z(n5187) );
  MUX2_X1 U5241 ( .A(reg_mem[138]), .B(reg_mem[130]), .S(n6768), .Z(n5188) );
  MUX2_X1 U5242 ( .A(reg_mem[154]), .B(reg_mem[146]), .S(n6781), .Z(n5189) );
  MUX2_X1 U5243 ( .A(n5189), .B(n5188), .S(n6723), .Z(n5190) );
  MUX2_X1 U5244 ( .A(reg_mem[170]), .B(reg_mem[162]), .S(n6775), .Z(n5191) );
  MUX2_X1 U5245 ( .A(reg_mem[186]), .B(reg_mem[178]), .S(n6774), .Z(n5192) );
  MUX2_X1 U5246 ( .A(n5192), .B(n5191), .S(n6719), .Z(n5193) );
  MUX2_X1 U5247 ( .A(n5193), .B(n5190), .S(n6717), .Z(n5194) );
  MUX2_X1 U5248 ( .A(reg_mem[202]), .B(reg_mem[194]), .S(n6746), .Z(n5195) );
  MUX2_X1 U5249 ( .A(reg_mem[218]), .B(reg_mem[210]), .S(n6747), .Z(n5196) );
  MUX2_X1 U5250 ( .A(n5196), .B(n5195), .S(n6720), .Z(n5197) );
  MUX2_X1 U5251 ( .A(reg_mem[234]), .B(reg_mem[226]), .S(n6749), .Z(n5198) );
  MUX2_X1 U5252 ( .A(reg_mem[250]), .B(reg_mem[242]), .S(n6772), .Z(n5199) );
  MUX2_X1 U5253 ( .A(n5199), .B(n5198), .S(n6739), .Z(n5200) );
  MUX2_X1 U5254 ( .A(n5200), .B(n5197), .S(n6717), .Z(n5201) );
  MUX2_X1 U5255 ( .A(n5201), .B(n5194), .S(n6704), .Z(n5202) );
  MUX2_X1 U5256 ( .A(n5202), .B(n5187), .S(n6700), .Z(n5203) );
  MUX2_X1 U5257 ( .A(reg_mem[266]), .B(reg_mem[258]), .S(n6769), .Z(n5204) );
  MUX2_X1 U5258 ( .A(reg_mem[282]), .B(reg_mem[274]), .S(n6744), .Z(n5205) );
  MUX2_X1 U5259 ( .A(n5205), .B(n5204), .S(n6724), .Z(n5206) );
  MUX2_X1 U5260 ( .A(reg_mem[298]), .B(reg_mem[290]), .S(n6764), .Z(n5207) );
  MUX2_X1 U5261 ( .A(reg_mem[314]), .B(reg_mem[306]), .S(n6749), .Z(n5208) );
  MUX2_X1 U5262 ( .A(n5208), .B(n5207), .S(n6719), .Z(n5209) );
  MUX2_X1 U5263 ( .A(n5209), .B(n5206), .S(n6717), .Z(n5210) );
  MUX2_X1 U5264 ( .A(reg_mem[330]), .B(reg_mem[322]), .S(n6770), .Z(n5211) );
  MUX2_X1 U5265 ( .A(reg_mem[346]), .B(reg_mem[338]), .S(n6748), .Z(n5212) );
  MUX2_X1 U5266 ( .A(n5212), .B(n5211), .S(n6718), .Z(n5213) );
  MUX2_X1 U5267 ( .A(reg_mem[362]), .B(reg_mem[354]), .S(n6764), .Z(n5214) );
  MUX2_X1 U5268 ( .A(reg_mem[378]), .B(reg_mem[370]), .S(n6766), .Z(n5215) );
  MUX2_X1 U5269 ( .A(n5215), .B(n5214), .S(addr_r[1]), .Z(n5216) );
  MUX2_X1 U5270 ( .A(n5216), .B(n5213), .S(n6717), .Z(n5217) );
  MUX2_X1 U5271 ( .A(n5217), .B(n5210), .S(n6703), .Z(n5218) );
  MUX2_X1 U5272 ( .A(reg_mem[394]), .B(reg_mem[386]), .S(n6779), .Z(n5219) );
  MUX2_X1 U5273 ( .A(reg_mem[410]), .B(reg_mem[402]), .S(n6768), .Z(n5220) );
  MUX2_X1 U5274 ( .A(n5220), .B(n5219), .S(n6721), .Z(n5221) );
  MUX2_X1 U5275 ( .A(reg_mem[426]), .B(reg_mem[418]), .S(n6767), .Z(n5222) );
  MUX2_X1 U5276 ( .A(reg_mem[442]), .B(reg_mem[434]), .S(n6755), .Z(n5223) );
  MUX2_X1 U5277 ( .A(n5223), .B(n5222), .S(n6735), .Z(n5224) );
  MUX2_X1 U5278 ( .A(n5224), .B(n5221), .S(n6717), .Z(n5225) );
  MUX2_X1 U5279 ( .A(reg_mem[458]), .B(reg_mem[450]), .S(n6762), .Z(n5226) );
  MUX2_X1 U5280 ( .A(reg_mem[474]), .B(reg_mem[466]), .S(n6745), .Z(n5227) );
  MUX2_X1 U5281 ( .A(n5227), .B(n5226), .S(n6736), .Z(n5228) );
  MUX2_X1 U5282 ( .A(reg_mem[490]), .B(reg_mem[482]), .S(n6754), .Z(n5229) );
  MUX2_X1 U5283 ( .A(reg_mem[506]), .B(reg_mem[498]), .S(n6767), .Z(n5230) );
  MUX2_X1 U5284 ( .A(n5230), .B(n5229), .S(n6725), .Z(n5231) );
  MUX2_X1 U5285 ( .A(n5231), .B(n5228), .S(n6717), .Z(n5232) );
  MUX2_X1 U5286 ( .A(n5232), .B(n5225), .S(n6705), .Z(n5233) );
  MUX2_X1 U5287 ( .A(n5233), .B(n5218), .S(n6700), .Z(n5234) );
  MUX2_X1 U5288 ( .A(n5234), .B(n5203), .S(n6697), .Z(n5235) );
  MUX2_X1 U5289 ( .A(reg_mem[522]), .B(reg_mem[514]), .S(n6777), .Z(n5236) );
  MUX2_X1 U5290 ( .A(reg_mem[538]), .B(reg_mem[530]), .S(n6743), .Z(n5237) );
  MUX2_X1 U5291 ( .A(n5237), .B(n5236), .S(n6736), .Z(n5238) );
  MUX2_X1 U5292 ( .A(reg_mem[554]), .B(reg_mem[546]), .S(n6765), .Z(n5239) );
  MUX2_X1 U5293 ( .A(reg_mem[570]), .B(reg_mem[562]), .S(n6753), .Z(n5240) );
  MUX2_X1 U5294 ( .A(n5240), .B(n5239), .S(n6727), .Z(n5241) );
  MUX2_X1 U5295 ( .A(n5241), .B(n5238), .S(n6707), .Z(n5242) );
  MUX2_X1 U5296 ( .A(reg_mem[586]), .B(reg_mem[578]), .S(n6775), .Z(n5243) );
  MUX2_X1 U5297 ( .A(reg_mem[602]), .B(reg_mem[594]), .S(n6782), .Z(n5244) );
  MUX2_X1 U5298 ( .A(n5244), .B(n5243), .S(n6721), .Z(n5245) );
  MUX2_X1 U5299 ( .A(reg_mem[618]), .B(reg_mem[610]), .S(n6752), .Z(n5246) );
  MUX2_X1 U5300 ( .A(reg_mem[634]), .B(reg_mem[626]), .S(n6757), .Z(n5247) );
  MUX2_X1 U5301 ( .A(n5247), .B(n5246), .S(n6718), .Z(n5248) );
  MUX2_X1 U5302 ( .A(n5248), .B(n5245), .S(n6708), .Z(n5249) );
  MUX2_X1 U5303 ( .A(n5249), .B(n5242), .S(addr_r[3]), .Z(n5250) );
  MUX2_X1 U5304 ( .A(reg_mem[650]), .B(reg_mem[642]), .S(n6750), .Z(n5251) );
  MUX2_X1 U5305 ( .A(reg_mem[666]), .B(reg_mem[658]), .S(n6743), .Z(n5252) );
  MUX2_X1 U5306 ( .A(n5252), .B(n5251), .S(n6734), .Z(n5253) );
  MUX2_X1 U5307 ( .A(reg_mem[682]), .B(reg_mem[674]), .S(n6779), .Z(n5254) );
  MUX2_X1 U5308 ( .A(reg_mem[698]), .B(reg_mem[690]), .S(n6760), .Z(n5255) );
  MUX2_X1 U5309 ( .A(n5255), .B(n5254), .S(n6733), .Z(n5256) );
  MUX2_X1 U5310 ( .A(n5256), .B(n5253), .S(n6717), .Z(n5257) );
  MUX2_X1 U5311 ( .A(reg_mem[714]), .B(reg_mem[706]), .S(n6782), .Z(n5258) );
  MUX2_X1 U5312 ( .A(reg_mem[730]), .B(reg_mem[722]), .S(n6762), .Z(n5259) );
  MUX2_X1 U5313 ( .A(n5259), .B(n5258), .S(n6722), .Z(n5260) );
  MUX2_X1 U5314 ( .A(reg_mem[746]), .B(reg_mem[738]), .S(n6745), .Z(n5261) );
  MUX2_X1 U5315 ( .A(reg_mem[762]), .B(reg_mem[754]), .S(n6759), .Z(n5262) );
  MUX2_X1 U5316 ( .A(n5262), .B(n5261), .S(n6734), .Z(n5263) );
  MUX2_X1 U5317 ( .A(n5263), .B(n5260), .S(n6711), .Z(n5264) );
  MUX2_X1 U5318 ( .A(n5264), .B(n5257), .S(n6701), .Z(n5265) );
  MUX2_X1 U5319 ( .A(n5265), .B(n5250), .S(addr_r[4]), .Z(n5266) );
  MUX2_X1 U5320 ( .A(reg_mem[778]), .B(reg_mem[770]), .S(n6768), .Z(n5267) );
  MUX2_X1 U5321 ( .A(reg_mem[794]), .B(reg_mem[786]), .S(n6754), .Z(n5268) );
  MUX2_X1 U5322 ( .A(n5268), .B(n5267), .S(n6723), .Z(n5269) );
  MUX2_X1 U5323 ( .A(reg_mem[810]), .B(reg_mem[802]), .S(n6760), .Z(n5270) );
  MUX2_X1 U5324 ( .A(reg_mem[826]), .B(reg_mem[818]), .S(n6777), .Z(n5271) );
  MUX2_X1 U5325 ( .A(n5271), .B(n5270), .S(n6723), .Z(n5272) );
  MUX2_X1 U5326 ( .A(n5272), .B(n5269), .S(addr_r[2]), .Z(n5273) );
  MUX2_X1 U5327 ( .A(reg_mem[842]), .B(reg_mem[834]), .S(n6773), .Z(n5274) );
  MUX2_X1 U5328 ( .A(reg_mem[858]), .B(reg_mem[850]), .S(n6769), .Z(n5275) );
  MUX2_X1 U5329 ( .A(n5275), .B(n5274), .S(n6739), .Z(n5276) );
  MUX2_X1 U5330 ( .A(reg_mem[874]), .B(reg_mem[866]), .S(n6779), .Z(n5277) );
  MUX2_X1 U5331 ( .A(reg_mem[890]), .B(reg_mem[882]), .S(n6744), .Z(n5278) );
  MUX2_X1 U5332 ( .A(n5278), .B(n5277), .S(n6722), .Z(n5279) );
  MUX2_X1 U5333 ( .A(n5279), .B(n5276), .S(n6710), .Z(n5280) );
  MUX2_X1 U5334 ( .A(n5280), .B(n5273), .S(n6706), .Z(n5281) );
  MUX2_X1 U5335 ( .A(reg_mem[906]), .B(reg_mem[898]), .S(n6781), .Z(n5282) );
  MUX2_X1 U5336 ( .A(reg_mem[922]), .B(reg_mem[914]), .S(n6768), .Z(n5283) );
  MUX2_X1 U5337 ( .A(n5283), .B(n5282), .S(n6739), .Z(n5284) );
  MUX2_X1 U5338 ( .A(reg_mem[938]), .B(reg_mem[930]), .S(n6771), .Z(n5285) );
  MUX2_X1 U5339 ( .A(reg_mem[954]), .B(reg_mem[946]), .S(n6781), .Z(n5286) );
  MUX2_X1 U5340 ( .A(n5286), .B(n5285), .S(n6739), .Z(n5287) );
  MUX2_X1 U5341 ( .A(n5287), .B(n5284), .S(n6709), .Z(n5288) );
  MUX2_X1 U5342 ( .A(reg_mem[970]), .B(reg_mem[962]), .S(n6746), .Z(n5289) );
  MUX2_X1 U5343 ( .A(reg_mem[986]), .B(reg_mem[978]), .S(n6770), .Z(n5290) );
  MUX2_X1 U5344 ( .A(n5290), .B(n5289), .S(n6727), .Z(n5291) );
  MUX2_X1 U5345 ( .A(reg_mem[1002]), .B(reg_mem[994]), .S(n6782), .Z(n5292) );
  MUX2_X1 U5346 ( .A(reg_mem[1018]), .B(reg_mem[1010]), .S(n6772), .Z(n5293)
         );
  MUX2_X1 U5347 ( .A(n5293), .B(n5292), .S(n6718), .Z(n5294) );
  MUX2_X1 U5348 ( .A(n5294), .B(n5291), .S(n6715), .Z(n5295) );
  MUX2_X1 U5349 ( .A(n5295), .B(n5288), .S(n6701), .Z(n5296) );
  MUX2_X1 U5350 ( .A(n5296), .B(n5281), .S(n6700), .Z(n5297) );
  MUX2_X1 U5351 ( .A(n5297), .B(n5266), .S(n6697), .Z(n5298) );
  MUX2_X1 U5352 ( .A(n5298), .B(n5235), .S(addr_r[6]), .Z(n5299) );
  MUX2_X1 U5353 ( .A(reg_mem[1034]), .B(reg_mem[1026]), .S(n6775), .Z(n5300)
         );
  MUX2_X1 U5354 ( .A(reg_mem[1050]), .B(reg_mem[1042]), .S(n6751), .Z(n5301)
         );
  MUX2_X1 U5355 ( .A(n5301), .B(n5300), .S(n6720), .Z(n5302) );
  MUX2_X1 U5356 ( .A(reg_mem[1066]), .B(reg_mem[1058]), .S(n6745), .Z(n5303)
         );
  MUX2_X1 U5357 ( .A(reg_mem[1082]), .B(reg_mem[1074]), .S(n6748), .Z(n5304)
         );
  MUX2_X1 U5358 ( .A(n5304), .B(n5303), .S(n6719), .Z(n5305) );
  MUX2_X1 U5359 ( .A(n5305), .B(n5302), .S(n6717), .Z(n5306) );
  MUX2_X1 U5360 ( .A(reg_mem[1098]), .B(reg_mem[1090]), .S(n6743), .Z(n5307)
         );
  MUX2_X1 U5361 ( .A(reg_mem[1114]), .B(reg_mem[1106]), .S(n6764), .Z(n5308)
         );
  MUX2_X1 U5362 ( .A(n5308), .B(n5307), .S(n6730), .Z(n5309) );
  MUX2_X1 U5363 ( .A(reg_mem[1130]), .B(reg_mem[1122]), .S(n6749), .Z(n5310)
         );
  MUX2_X1 U5364 ( .A(reg_mem[1146]), .B(reg_mem[1138]), .S(n6744), .Z(n5311)
         );
  MUX2_X1 U5365 ( .A(n5311), .B(n5310), .S(n6719), .Z(n5312) );
  MUX2_X1 U5366 ( .A(n5312), .B(n5309), .S(n6717), .Z(n5313) );
  MUX2_X1 U5367 ( .A(n5313), .B(n5306), .S(n6702), .Z(n5314) );
  MUX2_X1 U5368 ( .A(reg_mem[1162]), .B(reg_mem[1154]), .S(n6761), .Z(n5315)
         );
  MUX2_X1 U5369 ( .A(reg_mem[1178]), .B(reg_mem[1170]), .S(n6756), .Z(n5316)
         );
  MUX2_X1 U5370 ( .A(n5316), .B(n5315), .S(n6727), .Z(n5317) );
  MUX2_X1 U5371 ( .A(reg_mem[1194]), .B(reg_mem[1186]), .S(n6760), .Z(n5318)
         );
  MUX2_X1 U5372 ( .A(reg_mem[1210]), .B(reg_mem[1202]), .S(n6780), .Z(n5319)
         );
  MUX2_X1 U5373 ( .A(n5319), .B(n5318), .S(n6725), .Z(n5320) );
  MUX2_X1 U5374 ( .A(n5320), .B(n5317), .S(n6715), .Z(n5321) );
  MUX2_X1 U5375 ( .A(reg_mem[1226]), .B(reg_mem[1218]), .S(n6755), .Z(n5322)
         );
  MUX2_X1 U5376 ( .A(reg_mem[1242]), .B(reg_mem[1234]), .S(n6754), .Z(n5323)
         );
  MUX2_X1 U5377 ( .A(n5323), .B(n5322), .S(n6725), .Z(n5324) );
  MUX2_X1 U5378 ( .A(reg_mem[1258]), .B(reg_mem[1250]), .S(n6766), .Z(n5325)
         );
  MUX2_X1 U5379 ( .A(reg_mem[1274]), .B(reg_mem[1266]), .S(n6765), .Z(n5326)
         );
  MUX2_X1 U5380 ( .A(n5326), .B(n5325), .S(n6738), .Z(n5327) );
  MUX2_X1 U5381 ( .A(n5327), .B(n5324), .S(n6717), .Z(n5328) );
  MUX2_X1 U5382 ( .A(n5328), .B(n5321), .S(n6704), .Z(n5329) );
  MUX2_X1 U5383 ( .A(n5329), .B(n5314), .S(n6700), .Z(n5330) );
  MUX2_X1 U5384 ( .A(reg_mem[1290]), .B(reg_mem[1282]), .S(n6759), .Z(n5331)
         );
  MUX2_X1 U5385 ( .A(reg_mem[1306]), .B(reg_mem[1298]), .S(n6757), .Z(n5332)
         );
  MUX2_X1 U5386 ( .A(n5332), .B(n5331), .S(n6725), .Z(n5333) );
  MUX2_X1 U5387 ( .A(reg_mem[1322]), .B(reg_mem[1314]), .S(n6758), .Z(n5334)
         );
  MUX2_X1 U5388 ( .A(reg_mem[1338]), .B(reg_mem[1330]), .S(n6753), .Z(n5335)
         );
  MUX2_X1 U5389 ( .A(n5335), .B(n5334), .S(n6739), .Z(n5336) );
  MUX2_X1 U5390 ( .A(n5336), .B(n5333), .S(n6708), .Z(n5337) );
  MUX2_X1 U5391 ( .A(reg_mem[1354]), .B(reg_mem[1346]), .S(n6766), .Z(n5338)
         );
  MUX2_X1 U5392 ( .A(reg_mem[1370]), .B(reg_mem[1362]), .S(n6763), .Z(n5339)
         );
  MUX2_X1 U5393 ( .A(n5339), .B(n5338), .S(n6721), .Z(n5340) );
  MUX2_X1 U5394 ( .A(reg_mem[1386]), .B(reg_mem[1378]), .S(n6767), .Z(n5341)
         );
  MUX2_X1 U5395 ( .A(reg_mem[1402]), .B(reg_mem[1394]), .S(n6775), .Z(n5342)
         );
  MUX2_X1 U5396 ( .A(n5342), .B(n5341), .S(addr_r[1]), .Z(n5343) );
  MUX2_X1 U5397 ( .A(n5343), .B(n5340), .S(n6712), .Z(n5344) );
  MUX2_X1 U5398 ( .A(n5344), .B(n5337), .S(n6706), .Z(n5345) );
  MUX2_X1 U5399 ( .A(reg_mem[1418]), .B(reg_mem[1410]), .S(n6771), .Z(n5346)
         );
  MUX2_X1 U5400 ( .A(reg_mem[1434]), .B(reg_mem[1426]), .S(n6764), .Z(n5347)
         );
  MUX2_X1 U5401 ( .A(n5347), .B(n5346), .S(n6721), .Z(n5348) );
  MUX2_X1 U5402 ( .A(reg_mem[1450]), .B(reg_mem[1442]), .S(n6772), .Z(n5349)
         );
  MUX2_X1 U5403 ( .A(reg_mem[1466]), .B(reg_mem[1458]), .S(n6749), .Z(n5350)
         );
  MUX2_X1 U5404 ( .A(n5350), .B(n5349), .S(n6720), .Z(n5351) );
  MUX2_X1 U5405 ( .A(n5351), .B(n5348), .S(n6707), .Z(n5352) );
  MUX2_X1 U5406 ( .A(reg_mem[1482]), .B(reg_mem[1474]), .S(n6770), .Z(n5353)
         );
  MUX2_X1 U5407 ( .A(reg_mem[1498]), .B(reg_mem[1490]), .S(n6773), .Z(n5354)
         );
  MUX2_X1 U5408 ( .A(n5354), .B(n5353), .S(n6734), .Z(n5355) );
  MUX2_X1 U5409 ( .A(reg_mem[1514]), .B(reg_mem[1506]), .S(n6774), .Z(n5356)
         );
  MUX2_X1 U5410 ( .A(reg_mem[1530]), .B(reg_mem[1522]), .S(n6750), .Z(n5357)
         );
  MUX2_X1 U5411 ( .A(n5357), .B(n5356), .S(n6721), .Z(n5358) );
  MUX2_X1 U5412 ( .A(n5358), .B(n5355), .S(n6715), .Z(n5359) );
  MUX2_X1 U5413 ( .A(n5359), .B(n5352), .S(addr_r[3]), .Z(n5360) );
  MUX2_X1 U5414 ( .A(n5360), .B(n5345), .S(n6700), .Z(n5361) );
  MUX2_X1 U5415 ( .A(n5361), .B(n5330), .S(n6697), .Z(n5362) );
  MUX2_X1 U5416 ( .A(reg_mem[1546]), .B(reg_mem[1538]), .S(n6753), .Z(n5363)
         );
  MUX2_X1 U5417 ( .A(reg_mem[1562]), .B(reg_mem[1554]), .S(n6770), .Z(n5364)
         );
  MUX2_X1 U5418 ( .A(n5364), .B(n5363), .S(n6719), .Z(n5365) );
  MUX2_X1 U5419 ( .A(reg_mem[1578]), .B(reg_mem[1570]), .S(n6753), .Z(n5366)
         );
  MUX2_X1 U5420 ( .A(reg_mem[1594]), .B(reg_mem[1586]), .S(n6753), .Z(n5367)
         );
  MUX2_X1 U5421 ( .A(n5367), .B(n5366), .S(n6733), .Z(n5368) );
  MUX2_X1 U5422 ( .A(n5368), .B(n5365), .S(n6709), .Z(n5369) );
  MUX2_X1 U5423 ( .A(reg_mem[1610]), .B(reg_mem[1602]), .S(n6767), .Z(n5370)
         );
  MUX2_X1 U5424 ( .A(reg_mem[1626]), .B(reg_mem[1618]), .S(n6772), .Z(n5371)
         );
  MUX2_X1 U5425 ( .A(n5371), .B(n5370), .S(n6735), .Z(n5372) );
  MUX2_X1 U5426 ( .A(reg_mem[1642]), .B(reg_mem[1634]), .S(n6766), .Z(n5373)
         );
  MUX2_X1 U5427 ( .A(reg_mem[1658]), .B(reg_mem[1650]), .S(n6758), .Z(n5374)
         );
  MUX2_X1 U5428 ( .A(n5374), .B(n5373), .S(n6731), .Z(n5375) );
  MUX2_X1 U5429 ( .A(n5375), .B(n5372), .S(n6712), .Z(n5376) );
  MUX2_X1 U5430 ( .A(n5376), .B(n5369), .S(n6704), .Z(n5377) );
  MUX2_X1 U5431 ( .A(reg_mem[1674]), .B(reg_mem[1666]), .S(n6764), .Z(n5378)
         );
  MUX2_X1 U5432 ( .A(reg_mem[1690]), .B(reg_mem[1682]), .S(n6753), .Z(n5379)
         );
  MUX2_X1 U5433 ( .A(n5379), .B(n5378), .S(n6719), .Z(n5380) );
  MUX2_X1 U5434 ( .A(reg_mem[1706]), .B(reg_mem[1698]), .S(n6753), .Z(n5381)
         );
  MUX2_X1 U5435 ( .A(reg_mem[1722]), .B(reg_mem[1714]), .S(n6753), .Z(n5382)
         );
  MUX2_X1 U5436 ( .A(n5382), .B(n5381), .S(n6718), .Z(n5383) );
  MUX2_X1 U5437 ( .A(n5383), .B(n5380), .S(n6713), .Z(n5384) );
  MUX2_X1 U5438 ( .A(reg_mem[1738]), .B(reg_mem[1730]), .S(n6766), .Z(n5385)
         );
  MUX2_X1 U5439 ( .A(reg_mem[1754]), .B(reg_mem[1746]), .S(n6774), .Z(n5386)
         );
  MUX2_X1 U5440 ( .A(n5386), .B(n5385), .S(n6733), .Z(n5387) );
  MUX2_X1 U5441 ( .A(reg_mem[1770]), .B(reg_mem[1762]), .S(n6777), .Z(n5388)
         );
  MUX2_X1 U5442 ( .A(reg_mem[1786]), .B(reg_mem[1778]), .S(n6780), .Z(n5389)
         );
  MUX2_X1 U5443 ( .A(n5389), .B(n5388), .S(n6732), .Z(n5390) );
  MUX2_X1 U5444 ( .A(n5390), .B(n5387), .S(n6716), .Z(n5391) );
  MUX2_X1 U5445 ( .A(n5391), .B(n5384), .S(n6705), .Z(n5392) );
  MUX2_X1 U5446 ( .A(n5392), .B(n5377), .S(n6700), .Z(n5393) );
  MUX2_X1 U5447 ( .A(reg_mem[1802]), .B(reg_mem[1794]), .S(n6743), .Z(n5394)
         );
  MUX2_X1 U5448 ( .A(reg_mem[1818]), .B(reg_mem[1810]), .S(n6764), .Z(n5395)
         );
  MUX2_X1 U5449 ( .A(n5395), .B(n5394), .S(n6726), .Z(n5396) );
  MUX2_X1 U5450 ( .A(reg_mem[1834]), .B(reg_mem[1826]), .S(n6765), .Z(n5397)
         );
  MUX2_X1 U5451 ( .A(reg_mem[1850]), .B(reg_mem[1842]), .S(n6775), .Z(n5398)
         );
  MUX2_X1 U5452 ( .A(n5398), .B(n5397), .S(n6730), .Z(n5399) );
  MUX2_X1 U5453 ( .A(n5399), .B(n5396), .S(n6714), .Z(n5400) );
  MUX2_X1 U5454 ( .A(reg_mem[1866]), .B(reg_mem[1858]), .S(n6772), .Z(n5401)
         );
  MUX2_X1 U5455 ( .A(reg_mem[1882]), .B(reg_mem[1874]), .S(n6773), .Z(n5402)
         );
  MUX2_X1 U5456 ( .A(n5402), .B(n5401), .S(n6729), .Z(n5403) );
  MUX2_X1 U5457 ( .A(reg_mem[1898]), .B(reg_mem[1890]), .S(n6763), .Z(n5404)
         );
  MUX2_X1 U5458 ( .A(reg_mem[1914]), .B(reg_mem[1906]), .S(n6776), .Z(n5405)
         );
  MUX2_X1 U5459 ( .A(n5405), .B(n5404), .S(n6720), .Z(n5406) );
  MUX2_X1 U5460 ( .A(n5406), .B(n5403), .S(n6713), .Z(n5407) );
  MUX2_X1 U5461 ( .A(n5407), .B(n5400), .S(n6702), .Z(n5408) );
  MUX2_X1 U5462 ( .A(reg_mem[1930]), .B(reg_mem[1922]), .S(n6752), .Z(n5409)
         );
  MUX2_X1 U5463 ( .A(reg_mem[1946]), .B(reg_mem[1938]), .S(n6757), .Z(n5410)
         );
  MUX2_X1 U5464 ( .A(n5410), .B(n5409), .S(n6739), .Z(n5411) );
  MUX2_X1 U5465 ( .A(reg_mem[1962]), .B(reg_mem[1954]), .S(n6758), .Z(n5412)
         );
  MUX2_X1 U5466 ( .A(reg_mem[1978]), .B(reg_mem[1970]), .S(n6761), .Z(n5413)
         );
  MUX2_X1 U5467 ( .A(n5413), .B(n5412), .S(n6739), .Z(n5414) );
  MUX2_X1 U5468 ( .A(n5414), .B(n5411), .S(n6711), .Z(n5415) );
  MUX2_X1 U5469 ( .A(reg_mem[1994]), .B(reg_mem[1986]), .S(n6762), .Z(n5416)
         );
  MUX2_X1 U5470 ( .A(reg_mem[2010]), .B(reg_mem[2002]), .S(n6751), .Z(n5417)
         );
  MUX2_X1 U5471 ( .A(n5417), .B(n5416), .S(n6733), .Z(n5418) );
  MUX2_X1 U5472 ( .A(reg_mem[2026]), .B(reg_mem[2018]), .S(n6759), .Z(n5419)
         );
  MUX2_X1 U5473 ( .A(reg_mem[2042]), .B(reg_mem[2034]), .S(n6750), .Z(n5420)
         );
  MUX2_X1 U5474 ( .A(n5420), .B(n5419), .S(n6728), .Z(n5421) );
  MUX2_X1 U5475 ( .A(n5421), .B(n5418), .S(n6713), .Z(n5422) );
  MUX2_X1 U5476 ( .A(n5422), .B(n5415), .S(addr_r[3]), .Z(n5423) );
  MUX2_X1 U5477 ( .A(n5423), .B(n5408), .S(n6699), .Z(n5424) );
  MUX2_X1 U5478 ( .A(n5424), .B(n5393), .S(n6697), .Z(n5425) );
  MUX2_X1 U5479 ( .A(n5425), .B(n5362), .S(addr_r[6]), .Z(n5426) );
  MUX2_X1 U5480 ( .A(n5426), .B(n5299), .S(addr_r[7]), .Z(data_r[2]) );
  MUX2_X1 U5481 ( .A(reg_mem[11]), .B(reg_mem[3]), .S(n6743), .Z(n5427) );
  MUX2_X1 U5482 ( .A(reg_mem[27]), .B(reg_mem[19]), .S(n6778), .Z(n5428) );
  MUX2_X1 U5483 ( .A(n5428), .B(n5427), .S(n6734), .Z(n5429) );
  MUX2_X1 U5484 ( .A(reg_mem[43]), .B(reg_mem[35]), .S(n6781), .Z(n5430) );
  MUX2_X1 U5485 ( .A(reg_mem[59]), .B(reg_mem[51]), .S(n6782), .Z(n5431) );
  MUX2_X1 U5486 ( .A(n5431), .B(n5430), .S(n6729), .Z(n5432) );
  MUX2_X1 U5487 ( .A(n5432), .B(n5429), .S(n6711), .Z(n5433) );
  MUX2_X1 U5488 ( .A(reg_mem[75]), .B(reg_mem[67]), .S(n6754), .Z(n5434) );
  MUX2_X1 U5489 ( .A(reg_mem[91]), .B(reg_mem[83]), .S(n6762), .Z(n5435) );
  MUX2_X1 U5490 ( .A(n5435), .B(n5434), .S(n6718), .Z(n5436) );
  MUX2_X1 U5491 ( .A(reg_mem[107]), .B(reg_mem[99]), .S(n6757), .Z(n5437) );
  MUX2_X1 U5492 ( .A(reg_mem[123]), .B(reg_mem[115]), .S(n6761), .Z(n5438) );
  MUX2_X1 U5493 ( .A(n5438), .B(n5437), .S(n6732), .Z(n5439) );
  MUX2_X1 U5494 ( .A(n5439), .B(n5436), .S(n6707), .Z(n5440) );
  MUX2_X1 U5495 ( .A(n5440), .B(n5433), .S(n6703), .Z(n5441) );
  MUX2_X1 U5496 ( .A(reg_mem[139]), .B(reg_mem[131]), .S(n6761), .Z(n5442) );
  MUX2_X1 U5497 ( .A(reg_mem[155]), .B(reg_mem[147]), .S(n6756), .Z(n5443) );
  MUX2_X1 U5498 ( .A(n5443), .B(n5442), .S(n6732), .Z(n5444) );
  MUX2_X1 U5499 ( .A(reg_mem[171]), .B(reg_mem[163]), .S(n6760), .Z(n5445) );
  MUX2_X1 U5500 ( .A(reg_mem[187]), .B(reg_mem[179]), .S(n6758), .Z(n5446) );
  MUX2_X1 U5501 ( .A(n5446), .B(n5445), .S(n6734), .Z(n5447) );
  MUX2_X1 U5502 ( .A(n5447), .B(n5444), .S(n6711), .Z(n5448) );
  MUX2_X1 U5503 ( .A(reg_mem[203]), .B(reg_mem[195]), .S(n6752), .Z(n5449) );
  MUX2_X1 U5504 ( .A(reg_mem[219]), .B(reg_mem[211]), .S(n6751), .Z(n5450) );
  MUX2_X1 U5505 ( .A(n5450), .B(n5449), .S(n6720), .Z(n5451) );
  MUX2_X1 U5506 ( .A(reg_mem[235]), .B(reg_mem[227]), .S(n6759), .Z(n5452) );
  MUX2_X1 U5507 ( .A(reg_mem[251]), .B(reg_mem[243]), .S(n6750), .Z(n5453) );
  MUX2_X1 U5508 ( .A(n5453), .B(n5452), .S(n6739), .Z(n5454) );
  MUX2_X1 U5509 ( .A(n5454), .B(n5451), .S(n6709), .Z(n5455) );
  MUX2_X1 U5510 ( .A(n5455), .B(n5448), .S(n6706), .Z(n5456) );
  MUX2_X1 U5511 ( .A(n5456), .B(n5441), .S(n6699), .Z(n5457) );
  MUX2_X1 U5512 ( .A(reg_mem[267]), .B(reg_mem[259]), .S(n6761), .Z(n5458) );
  MUX2_X1 U5513 ( .A(reg_mem[283]), .B(reg_mem[275]), .S(n6744), .Z(n5459) );
  MUX2_X1 U5514 ( .A(n5459), .B(n5458), .S(n6721), .Z(n5460) );
  MUX2_X1 U5515 ( .A(reg_mem[299]), .B(reg_mem[291]), .S(n6770), .Z(n5461) );
  MUX2_X1 U5516 ( .A(reg_mem[315]), .B(reg_mem[307]), .S(n6747), .Z(n5462) );
  MUX2_X1 U5517 ( .A(n5462), .B(n5461), .S(n6733), .Z(n5463) );
  MUX2_X1 U5518 ( .A(n5463), .B(n5460), .S(n6707), .Z(n5464) );
  MUX2_X1 U5519 ( .A(reg_mem[331]), .B(reg_mem[323]), .S(n6772), .Z(n5465) );
  MUX2_X1 U5520 ( .A(reg_mem[347]), .B(reg_mem[339]), .S(n6747), .Z(n5466) );
  MUX2_X1 U5521 ( .A(n5466), .B(n5465), .S(n6722), .Z(n5467) );
  MUX2_X1 U5522 ( .A(reg_mem[363]), .B(reg_mem[355]), .S(n6772), .Z(n5468) );
  MUX2_X1 U5523 ( .A(reg_mem[379]), .B(reg_mem[371]), .S(n6763), .Z(n5469) );
  MUX2_X1 U5524 ( .A(n5469), .B(n5468), .S(n6732), .Z(n5470) );
  MUX2_X1 U5525 ( .A(n5470), .B(n5467), .S(n6712), .Z(n5471) );
  MUX2_X1 U5526 ( .A(n5471), .B(n5464), .S(n6702), .Z(n5472) );
  MUX2_X1 U5527 ( .A(reg_mem[395]), .B(reg_mem[387]), .S(n6746), .Z(n5473) );
  MUX2_X1 U5528 ( .A(reg_mem[411]), .B(reg_mem[403]), .S(n6743), .Z(n5474) );
  MUX2_X1 U5529 ( .A(n5474), .B(n5473), .S(n6735), .Z(n5475) );
  MUX2_X1 U5530 ( .A(reg_mem[427]), .B(reg_mem[419]), .S(n6745), .Z(n5476) );
  MUX2_X1 U5531 ( .A(reg_mem[443]), .B(reg_mem[435]), .S(n6752), .Z(n5477) );
  MUX2_X1 U5532 ( .A(n5477), .B(n5476), .S(n6721), .Z(n5478) );
  MUX2_X1 U5533 ( .A(n5478), .B(n5475), .S(n6716), .Z(n5479) );
  MUX2_X1 U5534 ( .A(reg_mem[459]), .B(reg_mem[451]), .S(n6769), .Z(n5480) );
  MUX2_X1 U5535 ( .A(reg_mem[475]), .B(reg_mem[467]), .S(n6750), .Z(n5481) );
  MUX2_X1 U5536 ( .A(n5481), .B(n5480), .S(n6728), .Z(n5482) );
  MUX2_X1 U5537 ( .A(reg_mem[491]), .B(reg_mem[483]), .S(n6754), .Z(n5483) );
  MUX2_X1 U5538 ( .A(reg_mem[507]), .B(reg_mem[499]), .S(n6776), .Z(n5484) );
  MUX2_X1 U5539 ( .A(n5484), .B(n5483), .S(n6720), .Z(n5485) );
  MUX2_X1 U5540 ( .A(n5485), .B(n5482), .S(n6715), .Z(n5486) );
  MUX2_X1 U5541 ( .A(n5486), .B(n5479), .S(n6703), .Z(n5487) );
  MUX2_X1 U5542 ( .A(n5487), .B(n5472), .S(n6699), .Z(n5488) );
  MUX2_X1 U5543 ( .A(n5488), .B(n5457), .S(n6697), .Z(n5489) );
  MUX2_X1 U5544 ( .A(reg_mem[523]), .B(reg_mem[515]), .S(n6753), .Z(n5490) );
  MUX2_X1 U5545 ( .A(reg_mem[539]), .B(reg_mem[531]), .S(n6782), .Z(n5491) );
  MUX2_X1 U5546 ( .A(n5491), .B(n5490), .S(n6718), .Z(n5492) );
  MUX2_X1 U5547 ( .A(reg_mem[555]), .B(reg_mem[547]), .S(n6757), .Z(n5493) );
  MUX2_X1 U5548 ( .A(reg_mem[571]), .B(reg_mem[563]), .S(n6774), .Z(n5494) );
  MUX2_X1 U5549 ( .A(n5494), .B(n5493), .S(n6731), .Z(n5495) );
  MUX2_X1 U5550 ( .A(n5495), .B(n5492), .S(n6716), .Z(n5496) );
  MUX2_X1 U5551 ( .A(reg_mem[587]), .B(reg_mem[579]), .S(n6755), .Z(n5497) );
  MUX2_X1 U5552 ( .A(reg_mem[603]), .B(reg_mem[595]), .S(n6751), .Z(n5498) );
  MUX2_X1 U5553 ( .A(n5498), .B(n5497), .S(n6735), .Z(n5499) );
  MUX2_X1 U5554 ( .A(reg_mem[619]), .B(reg_mem[611]), .S(n6749), .Z(n5500) );
  MUX2_X1 U5555 ( .A(reg_mem[635]), .B(reg_mem[627]), .S(n6766), .Z(n5501) );
  MUX2_X1 U5556 ( .A(n5501), .B(n5500), .S(n6739), .Z(n5502) );
  MUX2_X1 U5557 ( .A(n5502), .B(n5499), .S(n6712), .Z(n5503) );
  MUX2_X1 U5558 ( .A(n5503), .B(n5496), .S(n6702), .Z(n5504) );
  MUX2_X1 U5559 ( .A(reg_mem[651]), .B(reg_mem[643]), .S(n6757), .Z(n5505) );
  MUX2_X1 U5560 ( .A(reg_mem[667]), .B(reg_mem[659]), .S(n6777), .Z(n5506) );
  MUX2_X1 U5561 ( .A(n5506), .B(n5505), .S(n6720), .Z(n5507) );
  MUX2_X1 U5562 ( .A(reg_mem[683]), .B(reg_mem[675]), .S(n6744), .Z(n5508) );
  MUX2_X1 U5563 ( .A(reg_mem[699]), .B(reg_mem[691]), .S(n6765), .Z(n5509) );
  MUX2_X1 U5564 ( .A(n5509), .B(n5508), .S(n6735), .Z(n5510) );
  MUX2_X1 U5565 ( .A(n5510), .B(n5507), .S(n6710), .Z(n5511) );
  MUX2_X1 U5566 ( .A(reg_mem[715]), .B(reg_mem[707]), .S(n6778), .Z(n5512) );
  MUX2_X1 U5567 ( .A(reg_mem[731]), .B(reg_mem[723]), .S(n6777), .Z(n5513) );
  MUX2_X1 U5568 ( .A(n5513), .B(n5512), .S(n6739), .Z(n5514) );
  MUX2_X1 U5569 ( .A(reg_mem[747]), .B(reg_mem[739]), .S(n6778), .Z(n5515) );
  MUX2_X1 U5570 ( .A(reg_mem[763]), .B(reg_mem[755]), .S(n6772), .Z(n5516) );
  MUX2_X1 U5571 ( .A(n5516), .B(n5515), .S(n6739), .Z(n5517) );
  MUX2_X1 U5572 ( .A(n5517), .B(n5514), .S(n6711), .Z(n5518) );
  MUX2_X1 U5573 ( .A(n5518), .B(n5511), .S(n6705), .Z(n5519) );
  MUX2_X1 U5574 ( .A(n5519), .B(n5504), .S(addr_r[4]), .Z(n5520) );
  MUX2_X1 U5575 ( .A(reg_mem[779]), .B(reg_mem[771]), .S(n6743), .Z(n5521) );
  MUX2_X1 U5576 ( .A(reg_mem[795]), .B(reg_mem[787]), .S(n6746), .Z(n5522) );
  MUX2_X1 U5577 ( .A(n5522), .B(n5521), .S(n6720), .Z(n5523) );
  MUX2_X1 U5578 ( .A(reg_mem[811]), .B(reg_mem[803]), .S(n6751), .Z(n5524) );
  MUX2_X1 U5579 ( .A(reg_mem[827]), .B(reg_mem[819]), .S(n6751), .Z(n5525) );
  MUX2_X1 U5580 ( .A(n5525), .B(n5524), .S(n6727), .Z(n5526) );
  MUX2_X1 U5581 ( .A(n5526), .B(n5523), .S(n6712), .Z(n5527) );
  MUX2_X1 U5582 ( .A(reg_mem[843]), .B(reg_mem[835]), .S(n6755), .Z(n5528) );
  MUX2_X1 U5583 ( .A(reg_mem[859]), .B(reg_mem[851]), .S(n6751), .Z(n5529) );
  MUX2_X1 U5584 ( .A(n5529), .B(n5528), .S(n6730), .Z(n5530) );
  MUX2_X1 U5585 ( .A(reg_mem[875]), .B(reg_mem[867]), .S(n6766), .Z(n5531) );
  MUX2_X1 U5586 ( .A(reg_mem[891]), .B(reg_mem[883]), .S(n6745), .Z(n5532) );
  MUX2_X1 U5587 ( .A(n5532), .B(n5531), .S(n6734), .Z(n5533) );
  MUX2_X1 U5588 ( .A(n5533), .B(n5530), .S(n6713), .Z(n5534) );
  MUX2_X1 U5589 ( .A(n5534), .B(n5527), .S(n6706), .Z(n5535) );
  MUX2_X1 U5590 ( .A(reg_mem[907]), .B(reg_mem[899]), .S(n6778), .Z(n5536) );
  MUX2_X1 U5591 ( .A(reg_mem[923]), .B(reg_mem[915]), .S(n6743), .Z(n5537) );
  MUX2_X1 U5592 ( .A(n5537), .B(n5536), .S(n6721), .Z(n5538) );
  MUX2_X1 U5593 ( .A(reg_mem[939]), .B(reg_mem[931]), .S(n6765), .Z(n5539) );
  MUX2_X1 U5594 ( .A(reg_mem[955]), .B(reg_mem[947]), .S(n6748), .Z(n5540) );
  MUX2_X1 U5595 ( .A(n5540), .B(n5539), .S(n6732), .Z(n5541) );
  MUX2_X1 U5596 ( .A(n5541), .B(n5538), .S(n6710), .Z(n5542) );
  MUX2_X1 U5597 ( .A(reg_mem[971]), .B(reg_mem[963]), .S(n6763), .Z(n5543) );
  MUX2_X1 U5598 ( .A(reg_mem[987]), .B(reg_mem[979]), .S(n6747), .Z(n5544) );
  MUX2_X1 U5599 ( .A(n5544), .B(n5543), .S(n6731), .Z(n5545) );
  MUX2_X1 U5600 ( .A(reg_mem[1003]), .B(reg_mem[995]), .S(n6749), .Z(n5546) );
  MUX2_X1 U5601 ( .A(reg_mem[1019]), .B(reg_mem[1011]), .S(n6746), .Z(n5547)
         );
  MUX2_X1 U5602 ( .A(n5547), .B(n5546), .S(n6718), .Z(n5548) );
  MUX2_X1 U5603 ( .A(n5548), .B(n5545), .S(n6714), .Z(n5549) );
  MUX2_X1 U5604 ( .A(n5549), .B(n5542), .S(n6702), .Z(n5550) );
  MUX2_X1 U5605 ( .A(n5550), .B(n5535), .S(n6699), .Z(n5551) );
  MUX2_X1 U5606 ( .A(n5551), .B(n5520), .S(n6697), .Z(n5552) );
  MUX2_X1 U5607 ( .A(n5552), .B(n5489), .S(addr_r[6]), .Z(n5553) );
  MUX2_X1 U5608 ( .A(reg_mem[1035]), .B(reg_mem[1027]), .S(n6752), .Z(n5554)
         );
  MUX2_X1 U5609 ( .A(reg_mem[1051]), .B(reg_mem[1043]), .S(n6764), .Z(n5555)
         );
  MUX2_X1 U5610 ( .A(n5555), .B(n5554), .S(n6732), .Z(n5556) );
  MUX2_X1 U5611 ( .A(reg_mem[1067]), .B(reg_mem[1059]), .S(n6768), .Z(n5557)
         );
  MUX2_X1 U5612 ( .A(reg_mem[1083]), .B(reg_mem[1075]), .S(n6746), .Z(n5558)
         );
  MUX2_X1 U5613 ( .A(n5558), .B(n5557), .S(n6731), .Z(n5559) );
  MUX2_X1 U5614 ( .A(n5559), .B(n5556), .S(n6707), .Z(n5560) );
  MUX2_X1 U5615 ( .A(reg_mem[1099]), .B(reg_mem[1091]), .S(n6771), .Z(n5561)
         );
  MUX2_X1 U5616 ( .A(reg_mem[1115]), .B(reg_mem[1107]), .S(n6777), .Z(n5562)
         );
  MUX2_X1 U5617 ( .A(n5562), .B(n5561), .S(n6731), .Z(n5563) );
  MUX2_X1 U5618 ( .A(reg_mem[1131]), .B(reg_mem[1123]), .S(n6776), .Z(n5564)
         );
  MUX2_X1 U5619 ( .A(reg_mem[1147]), .B(reg_mem[1139]), .S(n6778), .Z(n5565)
         );
  MUX2_X1 U5620 ( .A(n5565), .B(n5564), .S(n6730), .Z(n5566) );
  MUX2_X1 U5621 ( .A(n5566), .B(n5563), .S(n6709), .Z(n5567) );
  MUX2_X1 U5622 ( .A(n5567), .B(n5560), .S(n6701), .Z(n5568) );
  MUX2_X1 U5623 ( .A(reg_mem[1163]), .B(reg_mem[1155]), .S(n6767), .Z(n5569)
         );
  MUX2_X1 U5624 ( .A(reg_mem[1179]), .B(reg_mem[1171]), .S(n6780), .Z(n5570)
         );
  MUX2_X1 U5625 ( .A(n5570), .B(n5569), .S(n6720), .Z(n5571) );
  MUX2_X1 U5626 ( .A(reg_mem[1195]), .B(reg_mem[1187]), .S(n6774), .Z(n5572)
         );
  MUX2_X1 U5627 ( .A(reg_mem[1211]), .B(reg_mem[1203]), .S(n6775), .Z(n5573)
         );
  MUX2_X1 U5628 ( .A(n5573), .B(n5572), .S(n6720), .Z(n5574) );
  MUX2_X1 U5629 ( .A(n5574), .B(n5571), .S(n6716), .Z(n5575) );
  MUX2_X1 U5630 ( .A(reg_mem[1227]), .B(reg_mem[1219]), .S(n6756), .Z(n5576)
         );
  MUX2_X1 U5631 ( .A(reg_mem[1243]), .B(reg_mem[1235]), .S(n6756), .Z(n5577)
         );
  MUX2_X1 U5632 ( .A(n5577), .B(n5576), .S(n6718), .Z(n5578) );
  MUX2_X1 U5633 ( .A(reg_mem[1259]), .B(reg_mem[1251]), .S(n6756), .Z(n5579)
         );
  MUX2_X1 U5634 ( .A(reg_mem[1275]), .B(reg_mem[1267]), .S(n6754), .Z(n5580)
         );
  MUX2_X1 U5635 ( .A(n5580), .B(n5579), .S(n6725), .Z(n5581) );
  MUX2_X1 U5636 ( .A(n5581), .B(n5578), .S(n6714), .Z(n5582) );
  MUX2_X1 U5637 ( .A(n5582), .B(n5575), .S(n6701), .Z(n5583) );
  MUX2_X1 U5638 ( .A(n5583), .B(n5568), .S(n6699), .Z(n5584) );
  MUX2_X1 U5639 ( .A(reg_mem[1291]), .B(reg_mem[1283]), .S(n6756), .Z(n5585)
         );
  MUX2_X1 U5640 ( .A(reg_mem[1307]), .B(reg_mem[1299]), .S(n6754), .Z(n5586)
         );
  MUX2_X1 U5641 ( .A(n5586), .B(n5585), .S(n6721), .Z(n5587) );
  MUX2_X1 U5642 ( .A(reg_mem[1323]), .B(reg_mem[1315]), .S(n6756), .Z(n5588)
         );
  MUX2_X1 U5643 ( .A(reg_mem[1339]), .B(reg_mem[1331]), .S(n6762), .Z(n5589)
         );
  MUX2_X1 U5644 ( .A(n5589), .B(n5588), .S(n6739), .Z(n5590) );
  MUX2_X1 U5645 ( .A(n5590), .B(n5587), .S(n6715), .Z(n5591) );
  MUX2_X1 U5646 ( .A(reg_mem[1355]), .B(reg_mem[1347]), .S(n6756), .Z(n5592)
         );
  MUX2_X1 U5647 ( .A(reg_mem[1371]), .B(reg_mem[1363]), .S(n6752), .Z(n5593)
         );
  MUX2_X1 U5648 ( .A(n5593), .B(n5592), .S(n6733), .Z(n5594) );
  MUX2_X1 U5649 ( .A(reg_mem[1387]), .B(reg_mem[1379]), .S(n6755), .Z(n5595)
         );
  MUX2_X1 U5650 ( .A(reg_mem[1403]), .B(reg_mem[1395]), .S(n6752), .Z(n5596)
         );
  MUX2_X1 U5651 ( .A(n5596), .B(n5595), .S(n6719), .Z(n5597) );
  MUX2_X1 U5652 ( .A(n5597), .B(n5594), .S(n6709), .Z(n5598) );
  MUX2_X1 U5653 ( .A(n5598), .B(n5591), .S(n6701), .Z(n5599) );
  MUX2_X1 U5654 ( .A(reg_mem[1419]), .B(reg_mem[1411]), .S(n6757), .Z(n5600)
         );
  MUX2_X1 U5655 ( .A(reg_mem[1435]), .B(reg_mem[1427]), .S(n6762), .Z(n5601)
         );
  MUX2_X1 U5656 ( .A(n5601), .B(n5600), .S(n6735), .Z(n5602) );
  MUX2_X1 U5657 ( .A(reg_mem[1451]), .B(reg_mem[1443]), .S(n6755), .Z(n5603)
         );
  MUX2_X1 U5658 ( .A(reg_mem[1467]), .B(reg_mem[1459]), .S(n6755), .Z(n5604)
         );
  MUX2_X1 U5659 ( .A(n5604), .B(n5603), .S(n6733), .Z(n5605) );
  MUX2_X1 U5660 ( .A(n5605), .B(n5602), .S(n6716), .Z(n5606) );
  MUX2_X1 U5661 ( .A(reg_mem[1483]), .B(reg_mem[1475]), .S(n6752), .Z(n5607)
         );
  MUX2_X1 U5662 ( .A(reg_mem[1499]), .B(reg_mem[1491]), .S(n6752), .Z(n5608)
         );
  MUX2_X1 U5663 ( .A(n5608), .B(n5607), .S(n6735), .Z(n5609) );
  MUX2_X1 U5664 ( .A(reg_mem[1515]), .B(reg_mem[1507]), .S(n6757), .Z(n5610)
         );
  MUX2_X1 U5665 ( .A(reg_mem[1531]), .B(reg_mem[1523]), .S(n6762), .Z(n5611)
         );
  MUX2_X1 U5666 ( .A(n5611), .B(n5610), .S(n6739), .Z(n5612) );
  MUX2_X1 U5667 ( .A(n5612), .B(n5609), .S(n6712), .Z(n5613) );
  MUX2_X1 U5668 ( .A(n5613), .B(n5606), .S(n6701), .Z(n5614) );
  MUX2_X1 U5669 ( .A(n5614), .B(n5599), .S(n6700), .Z(n5615) );
  MUX2_X1 U5670 ( .A(n5615), .B(n5584), .S(n6697), .Z(n5616) );
  MUX2_X1 U5671 ( .A(reg_mem[1547]), .B(reg_mem[1539]), .S(n6760), .Z(n5617)
         );
  MUX2_X1 U5672 ( .A(reg_mem[1563]), .B(reg_mem[1555]), .S(n6760), .Z(n5618)
         );
  MUX2_X1 U5673 ( .A(n5618), .B(n5617), .S(n6729), .Z(n5619) );
  MUX2_X1 U5674 ( .A(reg_mem[1579]), .B(reg_mem[1571]), .S(n6760), .Z(n5620)
         );
  MUX2_X1 U5675 ( .A(reg_mem[1595]), .B(reg_mem[1587]), .S(n6754), .Z(n5621)
         );
  MUX2_X1 U5676 ( .A(n5621), .B(n5620), .S(n6734), .Z(n5622) );
  MUX2_X1 U5677 ( .A(n5622), .B(n5619), .S(n6712), .Z(n5623) );
  MUX2_X1 U5678 ( .A(reg_mem[1611]), .B(reg_mem[1603]), .S(n6771), .Z(n5624)
         );
  MUX2_X1 U5679 ( .A(reg_mem[1627]), .B(reg_mem[1619]), .S(n6745), .Z(n5625)
         );
  MUX2_X1 U5680 ( .A(n5625), .B(n5624), .S(n6728), .Z(n5626) );
  MUX2_X1 U5681 ( .A(reg_mem[1643]), .B(reg_mem[1635]), .S(n6750), .Z(n5627)
         );
  MUX2_X1 U5682 ( .A(reg_mem[1659]), .B(reg_mem[1651]), .S(n6765), .Z(n5628)
         );
  MUX2_X1 U5683 ( .A(n5628), .B(n5627), .S(n6727), .Z(n5629) );
  MUX2_X1 U5684 ( .A(n5629), .B(n5626), .S(n6708), .Z(n5630) );
  MUX2_X1 U5685 ( .A(n5630), .B(n5623), .S(n6701), .Z(n5631) );
  MUX2_X1 U5686 ( .A(reg_mem[1675]), .B(reg_mem[1667]), .S(n6745), .Z(n5632)
         );
  MUX2_X1 U5687 ( .A(reg_mem[1691]), .B(reg_mem[1683]), .S(n6751), .Z(n5633)
         );
  MUX2_X1 U5688 ( .A(n5633), .B(n5632), .S(n6720), .Z(n5634) );
  MUX2_X1 U5689 ( .A(reg_mem[1707]), .B(reg_mem[1699]), .S(n6743), .Z(n5635)
         );
  MUX2_X1 U5690 ( .A(reg_mem[1723]), .B(reg_mem[1715]), .S(n6765), .Z(n5636)
         );
  MUX2_X1 U5691 ( .A(n5636), .B(n5635), .S(n6721), .Z(n5637) );
  MUX2_X1 U5692 ( .A(n5637), .B(n5634), .S(n6710), .Z(n5638) );
  MUX2_X1 U5693 ( .A(reg_mem[1739]), .B(reg_mem[1731]), .S(n6748), .Z(n5639)
         );
  MUX2_X1 U5694 ( .A(reg_mem[1755]), .B(reg_mem[1747]), .S(n6751), .Z(n5640)
         );
  MUX2_X1 U5695 ( .A(n5640), .B(n5639), .S(n6736), .Z(n5641) );
  MUX2_X1 U5696 ( .A(reg_mem[1771]), .B(reg_mem[1763]), .S(n6763), .Z(n5642)
         );
  MUX2_X1 U5697 ( .A(reg_mem[1787]), .B(reg_mem[1779]), .S(n6774), .Z(n5643)
         );
  MUX2_X1 U5698 ( .A(n5643), .B(n5642), .S(n6731), .Z(n5644) );
  MUX2_X1 U5699 ( .A(n5644), .B(n5641), .S(n6711), .Z(n5645) );
  MUX2_X1 U5700 ( .A(n5645), .B(n5638), .S(n6701), .Z(n5646) );
  MUX2_X1 U5701 ( .A(n5646), .B(n5631), .S(n6699), .Z(n5647) );
  MUX2_X1 U5702 ( .A(reg_mem[1803]), .B(reg_mem[1795]), .S(n6744), .Z(n5648)
         );
  MUX2_X1 U5703 ( .A(reg_mem[1819]), .B(reg_mem[1811]), .S(n6747), .Z(n5649)
         );
  MUX2_X1 U5704 ( .A(n5649), .B(n5648), .S(n6722), .Z(n5650) );
  MUX2_X1 U5705 ( .A(reg_mem[1835]), .B(reg_mem[1827]), .S(n6751), .Z(n5651)
         );
  MUX2_X1 U5706 ( .A(reg_mem[1851]), .B(reg_mem[1843]), .S(n6782), .Z(n5652)
         );
  MUX2_X1 U5707 ( .A(n5652), .B(n5651), .S(n6722), .Z(n5653) );
  MUX2_X1 U5708 ( .A(n5653), .B(n5650), .S(n6707), .Z(n5654) );
  MUX2_X1 U5709 ( .A(reg_mem[1867]), .B(reg_mem[1859]), .S(n6743), .Z(n5655)
         );
  MUX2_X1 U5710 ( .A(reg_mem[1883]), .B(reg_mem[1875]), .S(n6749), .Z(n5656)
         );
  MUX2_X1 U5711 ( .A(n5656), .B(n5655), .S(n6722), .Z(n5657) );
  MUX2_X1 U5712 ( .A(reg_mem[1899]), .B(reg_mem[1891]), .S(n6744), .Z(n5658)
         );
  MUX2_X1 U5713 ( .A(reg_mem[1915]), .B(reg_mem[1907]), .S(n6768), .Z(n5659)
         );
  MUX2_X1 U5714 ( .A(n5659), .B(n5658), .S(n6722), .Z(n5660) );
  MUX2_X1 U5715 ( .A(n5660), .B(n5657), .S(n6707), .Z(n5661) );
  MUX2_X1 U5716 ( .A(n5661), .B(n5654), .S(n6701), .Z(n5662) );
  MUX2_X1 U5717 ( .A(reg_mem[1931]), .B(reg_mem[1923]), .S(n6745), .Z(n5663)
         );
  MUX2_X1 U5718 ( .A(reg_mem[1947]), .B(reg_mem[1939]), .S(n6748), .Z(n5664)
         );
  MUX2_X1 U5719 ( .A(n5664), .B(n5663), .S(n6722), .Z(n5665) );
  MUX2_X1 U5720 ( .A(reg_mem[1963]), .B(reg_mem[1955]), .S(n6746), .Z(n5666)
         );
  MUX2_X1 U5721 ( .A(reg_mem[1979]), .B(reg_mem[1971]), .S(n6744), .Z(n5667)
         );
  MUX2_X1 U5722 ( .A(n5667), .B(n5666), .S(n6722), .Z(n5668) );
  MUX2_X1 U5723 ( .A(n5668), .B(n5665), .S(n6707), .Z(n5669) );
  MUX2_X1 U5724 ( .A(reg_mem[1995]), .B(reg_mem[1987]), .S(n6771), .Z(n5670)
         );
  MUX2_X1 U5725 ( .A(reg_mem[2011]), .B(reg_mem[2003]), .S(n6744), .Z(n5671)
         );
  MUX2_X1 U5726 ( .A(n5671), .B(n5670), .S(n6722), .Z(n5672) );
  MUX2_X1 U5727 ( .A(reg_mem[2027]), .B(reg_mem[2019]), .S(n6747), .Z(n5673)
         );
  MUX2_X1 U5728 ( .A(reg_mem[2043]), .B(reg_mem[2035]), .S(n6746), .Z(n5674)
         );
  MUX2_X1 U5729 ( .A(n5674), .B(n5673), .S(n6722), .Z(n5675) );
  MUX2_X1 U5730 ( .A(n5675), .B(n5672), .S(n6707), .Z(n5676) );
  MUX2_X1 U5731 ( .A(n5676), .B(n5669), .S(n6701), .Z(n5677) );
  MUX2_X1 U5732 ( .A(n5677), .B(n5662), .S(addr_r[4]), .Z(n5678) );
  MUX2_X1 U5733 ( .A(n5678), .B(n5647), .S(n6697), .Z(n5679) );
  MUX2_X1 U5734 ( .A(n5679), .B(n5616), .S(addr_r[6]), .Z(n5680) );
  MUX2_X1 U5735 ( .A(n5680), .B(n5553), .S(addr_r[7]), .Z(data_r[3]) );
  MUX2_X1 U5736 ( .A(reg_mem[12]), .B(reg_mem[4]), .S(n6762), .Z(n5681) );
  MUX2_X1 U5737 ( .A(reg_mem[28]), .B(reg_mem[20]), .S(n6757), .Z(n5682) );
  MUX2_X1 U5738 ( .A(n5682), .B(n5681), .S(n6722), .Z(n5683) );
  MUX2_X1 U5739 ( .A(reg_mem[44]), .B(reg_mem[36]), .S(n6755), .Z(n5684) );
  MUX2_X1 U5740 ( .A(reg_mem[60]), .B(reg_mem[52]), .S(n6752), .Z(n5685) );
  MUX2_X1 U5741 ( .A(n5685), .B(n5684), .S(n6722), .Z(n5686) );
  MUX2_X1 U5742 ( .A(n5686), .B(n5683), .S(n6707), .Z(n5687) );
  MUX2_X1 U5743 ( .A(reg_mem[76]), .B(reg_mem[68]), .S(n6752), .Z(n5688) );
  MUX2_X1 U5744 ( .A(reg_mem[92]), .B(reg_mem[84]), .S(n6754), .Z(n5689) );
  MUX2_X1 U5745 ( .A(n5689), .B(n5688), .S(n6722), .Z(n5690) );
  MUX2_X1 U5746 ( .A(reg_mem[108]), .B(reg_mem[100]), .S(n6755), .Z(n5691) );
  MUX2_X1 U5747 ( .A(reg_mem[124]), .B(reg_mem[116]), .S(n6757), .Z(n5692) );
  MUX2_X1 U5748 ( .A(n5692), .B(n5691), .S(n6722), .Z(n5693) );
  MUX2_X1 U5749 ( .A(n5693), .B(n5690), .S(n6707), .Z(n5694) );
  MUX2_X1 U5750 ( .A(n5694), .B(n5687), .S(n6701), .Z(n5695) );
  MUX2_X1 U5751 ( .A(reg_mem[140]), .B(reg_mem[132]), .S(n6776), .Z(n5696) );
  MUX2_X1 U5752 ( .A(reg_mem[156]), .B(reg_mem[148]), .S(n6777), .Z(n5697) );
  MUX2_X1 U5753 ( .A(n5697), .B(n5696), .S(n6737), .Z(n5698) );
  MUX2_X1 U5754 ( .A(reg_mem[172]), .B(reg_mem[164]), .S(n6781), .Z(n5699) );
  MUX2_X1 U5755 ( .A(reg_mem[188]), .B(reg_mem[180]), .S(n6773), .Z(n5700) );
  MUX2_X1 U5756 ( .A(n5700), .B(n5699), .S(n6736), .Z(n5701) );
  MUX2_X1 U5757 ( .A(n5701), .B(n5698), .S(n6707), .Z(n5702) );
  MUX2_X1 U5758 ( .A(reg_mem[204]), .B(reg_mem[196]), .S(n6779), .Z(n5703) );
  MUX2_X1 U5759 ( .A(reg_mem[220]), .B(reg_mem[212]), .S(n6770), .Z(n5704) );
  MUX2_X1 U5760 ( .A(n5704), .B(n5703), .S(n6730), .Z(n5705) );
  MUX2_X1 U5761 ( .A(reg_mem[236]), .B(reg_mem[228]), .S(n6766), .Z(n5706) );
  MUX2_X1 U5762 ( .A(reg_mem[252]), .B(reg_mem[244]), .S(n6767), .Z(n5707) );
  MUX2_X1 U5763 ( .A(n5707), .B(n5706), .S(n6727), .Z(n5708) );
  MUX2_X1 U5764 ( .A(n5708), .B(n5705), .S(n6707), .Z(n5709) );
  MUX2_X1 U5765 ( .A(n5709), .B(n5702), .S(n6701), .Z(n5710) );
  MUX2_X1 U5766 ( .A(n5710), .B(n5695), .S(n6699), .Z(n5711) );
  MUX2_X1 U5767 ( .A(reg_mem[268]), .B(reg_mem[260]), .S(n6771), .Z(n5712) );
  MUX2_X1 U5768 ( .A(reg_mem[284]), .B(reg_mem[276]), .S(n6778), .Z(n5713) );
  MUX2_X1 U5769 ( .A(n5713), .B(n5712), .S(n6736), .Z(n5714) );
  MUX2_X1 U5770 ( .A(reg_mem[300]), .B(reg_mem[292]), .S(n6782), .Z(n5715) );
  MUX2_X1 U5771 ( .A(reg_mem[316]), .B(reg_mem[308]), .S(n6763), .Z(n5716) );
  MUX2_X1 U5772 ( .A(n5716), .B(n5715), .S(n6738), .Z(n5717) );
  MUX2_X1 U5773 ( .A(n5717), .B(n5714), .S(n6707), .Z(n5718) );
  MUX2_X1 U5774 ( .A(reg_mem[332]), .B(reg_mem[324]), .S(n6743), .Z(n5719) );
  MUX2_X1 U5775 ( .A(reg_mem[348]), .B(reg_mem[340]), .S(n6743), .Z(n5720) );
  MUX2_X1 U5776 ( .A(n5720), .B(n5719), .S(n6728), .Z(n5721) );
  MUX2_X1 U5777 ( .A(reg_mem[364]), .B(reg_mem[356]), .S(n6743), .Z(n5722) );
  MUX2_X1 U5778 ( .A(reg_mem[380]), .B(reg_mem[372]), .S(n6743), .Z(n5723) );
  MUX2_X1 U5779 ( .A(n5723), .B(n5722), .S(n6726), .Z(n5724) );
  MUX2_X1 U5780 ( .A(n5724), .B(n5721), .S(n6707), .Z(n5725) );
  MUX2_X1 U5781 ( .A(n5725), .B(n5718), .S(n6701), .Z(n5726) );
  MUX2_X1 U5782 ( .A(reg_mem[396]), .B(reg_mem[388]), .S(n6743), .Z(n5727) );
  MUX2_X1 U5783 ( .A(reg_mem[412]), .B(reg_mem[404]), .S(n6743), .Z(n5728) );
  MUX2_X1 U5784 ( .A(n5728), .B(n5727), .S(n6729), .Z(n5729) );
  MUX2_X1 U5785 ( .A(reg_mem[428]), .B(reg_mem[420]), .S(n6743), .Z(n5730) );
  MUX2_X1 U5786 ( .A(reg_mem[444]), .B(reg_mem[436]), .S(n6743), .Z(n5731) );
  MUX2_X1 U5787 ( .A(n5731), .B(n5730), .S(n6728), .Z(n5732) );
  MUX2_X1 U5788 ( .A(n5732), .B(n5729), .S(n6707), .Z(n5733) );
  MUX2_X1 U5789 ( .A(reg_mem[460]), .B(reg_mem[452]), .S(n6743), .Z(n5734) );
  MUX2_X1 U5790 ( .A(reg_mem[476]), .B(reg_mem[468]), .S(n6743), .Z(n5735) );
  MUX2_X1 U5791 ( .A(n5735), .B(n5734), .S(n6737), .Z(n5736) );
  MUX2_X1 U5792 ( .A(reg_mem[492]), .B(reg_mem[484]), .S(n6743), .Z(n5737) );
  MUX2_X1 U5793 ( .A(reg_mem[508]), .B(reg_mem[500]), .S(n6743), .Z(n5738) );
  MUX2_X1 U5794 ( .A(n5738), .B(n5737), .S(n6719), .Z(n5739) );
  MUX2_X1 U5795 ( .A(n5739), .B(n5736), .S(n6707), .Z(n5740) );
  MUX2_X1 U5796 ( .A(n5740), .B(n5733), .S(n6701), .Z(n5741) );
  MUX2_X1 U5797 ( .A(n5741), .B(n5726), .S(n6699), .Z(n5742) );
  MUX2_X1 U5798 ( .A(n5742), .B(n5711), .S(n6697), .Z(n5743) );
  MUX2_X1 U5799 ( .A(reg_mem[524]), .B(reg_mem[516]), .S(n6744), .Z(n5744) );
  MUX2_X1 U5800 ( .A(reg_mem[540]), .B(reg_mem[532]), .S(n6744), .Z(n5745) );
  MUX2_X1 U5801 ( .A(n5745), .B(n5744), .S(n6723), .Z(n5746) );
  MUX2_X1 U5802 ( .A(reg_mem[556]), .B(reg_mem[548]), .S(n6744), .Z(n5747) );
  MUX2_X1 U5803 ( .A(reg_mem[572]), .B(reg_mem[564]), .S(n6744), .Z(n5748) );
  MUX2_X1 U5804 ( .A(n5748), .B(n5747), .S(n6723), .Z(n5749) );
  MUX2_X1 U5805 ( .A(n5749), .B(n5746), .S(n6708), .Z(n5750) );
  MUX2_X1 U5806 ( .A(reg_mem[588]), .B(reg_mem[580]), .S(n6744), .Z(n5751) );
  MUX2_X1 U5807 ( .A(reg_mem[604]), .B(reg_mem[596]), .S(n6744), .Z(n5752) );
  MUX2_X1 U5808 ( .A(n5752), .B(n5751), .S(n6723), .Z(n5753) );
  MUX2_X1 U5809 ( .A(reg_mem[620]), .B(reg_mem[612]), .S(n6744), .Z(n5754) );
  MUX2_X1 U5810 ( .A(reg_mem[636]), .B(reg_mem[628]), .S(n6744), .Z(n5755) );
  MUX2_X1 U5811 ( .A(n5755), .B(n5754), .S(n6723), .Z(n5756) );
  MUX2_X1 U5812 ( .A(n5756), .B(n5753), .S(n6708), .Z(n5757) );
  MUX2_X1 U5813 ( .A(n5757), .B(n5750), .S(n6702), .Z(n5758) );
  MUX2_X1 U5814 ( .A(reg_mem[652]), .B(reg_mem[644]), .S(n6744), .Z(n5759) );
  MUX2_X1 U5815 ( .A(reg_mem[668]), .B(reg_mem[660]), .S(n6744), .Z(n5760) );
  MUX2_X1 U5816 ( .A(n5760), .B(n5759), .S(n6723), .Z(n5761) );
  MUX2_X1 U5817 ( .A(reg_mem[684]), .B(reg_mem[676]), .S(n6744), .Z(n5762) );
  MUX2_X1 U5818 ( .A(reg_mem[700]), .B(reg_mem[692]), .S(n6744), .Z(n5763) );
  MUX2_X1 U5819 ( .A(n5763), .B(n5762), .S(n6723), .Z(n5764) );
  MUX2_X1 U5820 ( .A(n5764), .B(n5761), .S(n6708), .Z(n5765) );
  MUX2_X1 U5821 ( .A(reg_mem[716]), .B(reg_mem[708]), .S(n6745), .Z(n5766) );
  MUX2_X1 U5822 ( .A(reg_mem[732]), .B(reg_mem[724]), .S(n6745), .Z(n5767) );
  MUX2_X1 U5823 ( .A(n5767), .B(n5766), .S(n6723), .Z(n5768) );
  MUX2_X1 U5824 ( .A(reg_mem[748]), .B(reg_mem[740]), .S(n6745), .Z(n5769) );
  MUX2_X1 U5825 ( .A(reg_mem[764]), .B(reg_mem[756]), .S(n6745), .Z(n5770) );
  MUX2_X1 U5826 ( .A(n5770), .B(n5769), .S(n6723), .Z(n5771) );
  MUX2_X1 U5827 ( .A(n5771), .B(n5768), .S(n6708), .Z(n5772) );
  MUX2_X1 U5828 ( .A(n5772), .B(n5765), .S(n6702), .Z(n5773) );
  MUX2_X1 U5829 ( .A(n5773), .B(n5758), .S(n6699), .Z(n5774) );
  MUX2_X1 U5830 ( .A(reg_mem[780]), .B(reg_mem[772]), .S(n6745), .Z(n5775) );
  MUX2_X1 U5831 ( .A(reg_mem[796]), .B(reg_mem[788]), .S(n6745), .Z(n5776) );
  MUX2_X1 U5832 ( .A(n5776), .B(n5775), .S(n6723), .Z(n5777) );
  MUX2_X1 U5833 ( .A(reg_mem[812]), .B(reg_mem[804]), .S(n6745), .Z(n5778) );
  MUX2_X1 U5834 ( .A(reg_mem[828]), .B(reg_mem[820]), .S(n6745), .Z(n5779) );
  MUX2_X1 U5835 ( .A(n5779), .B(n5778), .S(n6723), .Z(n5780) );
  MUX2_X1 U5836 ( .A(n5780), .B(n5777), .S(n6708), .Z(n5781) );
  MUX2_X1 U5837 ( .A(reg_mem[844]), .B(reg_mem[836]), .S(n6745), .Z(n5782) );
  MUX2_X1 U5838 ( .A(reg_mem[860]), .B(reg_mem[852]), .S(n6745), .Z(n5783) );
  MUX2_X1 U5839 ( .A(n5783), .B(n5782), .S(n6723), .Z(n5784) );
  MUX2_X1 U5840 ( .A(reg_mem[876]), .B(reg_mem[868]), .S(n6745), .Z(n5785) );
  MUX2_X1 U5841 ( .A(reg_mem[892]), .B(reg_mem[884]), .S(n6745), .Z(n5786) );
  MUX2_X1 U5842 ( .A(n5786), .B(n5785), .S(n6723), .Z(n5787) );
  MUX2_X1 U5843 ( .A(n5787), .B(n5784), .S(n6708), .Z(n5788) );
  MUX2_X1 U5844 ( .A(n5788), .B(n5781), .S(n6702), .Z(n5789) );
  MUX2_X1 U5845 ( .A(reg_mem[908]), .B(reg_mem[900]), .S(n6746), .Z(n5790) );
  MUX2_X1 U5846 ( .A(reg_mem[924]), .B(reg_mem[916]), .S(n6746), .Z(n5791) );
  MUX2_X1 U5847 ( .A(n5791), .B(n5790), .S(n6724), .Z(n5792) );
  MUX2_X1 U5848 ( .A(reg_mem[940]), .B(reg_mem[932]), .S(n6746), .Z(n5793) );
  MUX2_X1 U5849 ( .A(reg_mem[956]), .B(reg_mem[948]), .S(n6746), .Z(n5794) );
  MUX2_X1 U5850 ( .A(n5794), .B(n5793), .S(n6724), .Z(n5795) );
  MUX2_X1 U5851 ( .A(n5795), .B(n5792), .S(n6708), .Z(n5796) );
  MUX2_X1 U5852 ( .A(reg_mem[972]), .B(reg_mem[964]), .S(n6746), .Z(n5797) );
  MUX2_X1 U5853 ( .A(reg_mem[988]), .B(reg_mem[980]), .S(n6746), .Z(n5798) );
  MUX2_X1 U5854 ( .A(n5798), .B(n5797), .S(n6724), .Z(n5799) );
  MUX2_X1 U5855 ( .A(reg_mem[1004]), .B(reg_mem[996]), .S(n6746), .Z(n5800) );
  MUX2_X1 U5856 ( .A(reg_mem[1020]), .B(reg_mem[1012]), .S(n6746), .Z(n5801)
         );
  MUX2_X1 U5857 ( .A(n5801), .B(n5800), .S(n6724), .Z(n5802) );
  MUX2_X1 U5858 ( .A(n5802), .B(n5799), .S(n6708), .Z(n5803) );
  MUX2_X1 U5859 ( .A(n5803), .B(n5796), .S(n6702), .Z(n5804) );
  MUX2_X1 U5860 ( .A(n5804), .B(n5789), .S(n6700), .Z(n5805) );
  MUX2_X1 U5861 ( .A(n5805), .B(n5774), .S(n6697), .Z(n5806) );
  MUX2_X1 U5862 ( .A(n5806), .B(n5743), .S(addr_r[6]), .Z(n5807) );
  MUX2_X1 U5863 ( .A(reg_mem[1036]), .B(reg_mem[1028]), .S(n6746), .Z(n5808)
         );
  MUX2_X1 U5864 ( .A(reg_mem[1052]), .B(reg_mem[1044]), .S(n6746), .Z(n5809)
         );
  MUX2_X1 U5865 ( .A(n5809), .B(n5808), .S(n6724), .Z(n5810) );
  MUX2_X1 U5866 ( .A(reg_mem[1068]), .B(reg_mem[1060]), .S(n6746), .Z(n5811)
         );
  MUX2_X1 U5867 ( .A(reg_mem[1084]), .B(reg_mem[1076]), .S(n6746), .Z(n5812)
         );
  MUX2_X1 U5868 ( .A(n5812), .B(n5811), .S(n6724), .Z(n5813) );
  MUX2_X1 U5869 ( .A(n5813), .B(n5810), .S(n6708), .Z(n5814) );
  MUX2_X1 U5870 ( .A(reg_mem[1100]), .B(reg_mem[1092]), .S(n6747), .Z(n5815)
         );
  MUX2_X1 U5871 ( .A(reg_mem[1116]), .B(reg_mem[1108]), .S(n6747), .Z(n5816)
         );
  MUX2_X1 U5872 ( .A(n5816), .B(n5815), .S(n6724), .Z(n5817) );
  MUX2_X1 U5873 ( .A(reg_mem[1132]), .B(reg_mem[1124]), .S(n6747), .Z(n5818)
         );
  MUX2_X1 U5874 ( .A(reg_mem[1148]), .B(reg_mem[1140]), .S(n6747), .Z(n5819)
         );
  MUX2_X1 U5875 ( .A(n5819), .B(n5818), .S(n6724), .Z(n5820) );
  MUX2_X1 U5876 ( .A(n5820), .B(n5817), .S(n6708), .Z(n5821) );
  MUX2_X1 U5877 ( .A(n5821), .B(n5814), .S(n6702), .Z(n5822) );
  MUX2_X1 U5878 ( .A(reg_mem[1164]), .B(reg_mem[1156]), .S(n6747), .Z(n5823)
         );
  MUX2_X1 U5879 ( .A(reg_mem[1180]), .B(reg_mem[1172]), .S(n6747), .Z(n5824)
         );
  MUX2_X1 U5880 ( .A(n5824), .B(n5823), .S(n6724), .Z(n5825) );
  MUX2_X1 U5881 ( .A(reg_mem[1196]), .B(reg_mem[1188]), .S(n6747), .Z(n5826)
         );
  MUX2_X1 U5882 ( .A(reg_mem[1212]), .B(reg_mem[1204]), .S(n6747), .Z(n5827)
         );
  MUX2_X1 U5883 ( .A(n5827), .B(n5826), .S(n6724), .Z(n5828) );
  MUX2_X1 U5884 ( .A(n5828), .B(n5825), .S(n6708), .Z(n5829) );
  MUX2_X1 U5885 ( .A(reg_mem[1228]), .B(reg_mem[1220]), .S(n6747), .Z(n5830)
         );
  MUX2_X1 U5886 ( .A(reg_mem[1244]), .B(reg_mem[1236]), .S(n6747), .Z(n5831)
         );
  MUX2_X1 U5887 ( .A(n5831), .B(n5830), .S(n6724), .Z(n5832) );
  MUX2_X1 U5888 ( .A(reg_mem[1260]), .B(reg_mem[1252]), .S(n6747), .Z(n5833)
         );
  MUX2_X1 U5889 ( .A(reg_mem[1276]), .B(reg_mem[1268]), .S(n6747), .Z(n5834)
         );
  MUX2_X1 U5890 ( .A(n5834), .B(n5833), .S(n6724), .Z(n5835) );
  MUX2_X1 U5891 ( .A(n5835), .B(n5832), .S(n6708), .Z(n5836) );
  MUX2_X1 U5892 ( .A(n5836), .B(n5829), .S(n6702), .Z(n5837) );
  MUX2_X1 U5893 ( .A(n5837), .B(n5822), .S(n6699), .Z(n5838) );
  MUX2_X1 U5894 ( .A(reg_mem[1292]), .B(reg_mem[1284]), .S(n6748), .Z(n5839)
         );
  MUX2_X1 U5895 ( .A(reg_mem[1308]), .B(reg_mem[1300]), .S(n6748), .Z(n5840)
         );
  MUX2_X1 U5896 ( .A(n5840), .B(n5839), .S(n6725), .Z(n5841) );
  MUX2_X1 U5897 ( .A(reg_mem[1324]), .B(reg_mem[1316]), .S(n6748), .Z(n5842)
         );
  MUX2_X1 U5898 ( .A(reg_mem[1340]), .B(reg_mem[1332]), .S(n6748), .Z(n5843)
         );
  MUX2_X1 U5899 ( .A(n5843), .B(n5842), .S(n6725), .Z(n5844) );
  MUX2_X1 U5900 ( .A(n5844), .B(n5841), .S(n6709), .Z(n5845) );
  MUX2_X1 U5901 ( .A(reg_mem[1356]), .B(reg_mem[1348]), .S(n6748), .Z(n5846)
         );
  MUX2_X1 U5902 ( .A(reg_mem[1372]), .B(reg_mem[1364]), .S(n6748), .Z(n5847)
         );
  MUX2_X1 U5903 ( .A(n5847), .B(n5846), .S(n6725), .Z(n5848) );
  MUX2_X1 U5904 ( .A(reg_mem[1388]), .B(reg_mem[1380]), .S(n6748), .Z(n5849)
         );
  MUX2_X1 U5905 ( .A(reg_mem[1404]), .B(reg_mem[1396]), .S(n6748), .Z(n5850)
         );
  MUX2_X1 U5906 ( .A(n5850), .B(n5849), .S(n6725), .Z(n5851) );
  MUX2_X1 U5907 ( .A(n5851), .B(n5848), .S(n6709), .Z(n5852) );
  MUX2_X1 U5908 ( .A(n5852), .B(n5845), .S(n6702), .Z(n5853) );
  MUX2_X1 U5909 ( .A(reg_mem[1420]), .B(reg_mem[1412]), .S(n6748), .Z(n5854)
         );
  MUX2_X1 U5910 ( .A(reg_mem[1436]), .B(reg_mem[1428]), .S(n6748), .Z(n5855)
         );
  MUX2_X1 U5911 ( .A(n5855), .B(n5854), .S(n6725), .Z(n5856) );
  MUX2_X1 U5912 ( .A(reg_mem[1452]), .B(reg_mem[1444]), .S(n6748), .Z(n5857)
         );
  MUX2_X1 U5913 ( .A(reg_mem[1468]), .B(reg_mem[1460]), .S(n6748), .Z(n5858)
         );
  MUX2_X1 U5914 ( .A(n5858), .B(n5857), .S(n6725), .Z(n5859) );
  MUX2_X1 U5915 ( .A(n5859), .B(n5856), .S(n6709), .Z(n5860) );
  MUX2_X1 U5916 ( .A(reg_mem[1484]), .B(reg_mem[1476]), .S(n6775), .Z(n5861)
         );
  MUX2_X1 U5917 ( .A(reg_mem[1500]), .B(reg_mem[1492]), .S(n6776), .Z(n5862)
         );
  MUX2_X1 U5918 ( .A(n5862), .B(n5861), .S(n6725), .Z(n5863) );
  MUX2_X1 U5919 ( .A(reg_mem[1516]), .B(reg_mem[1508]), .S(n6781), .Z(n5864)
         );
  MUX2_X1 U5920 ( .A(reg_mem[1532]), .B(reg_mem[1524]), .S(n6781), .Z(n5865)
         );
  MUX2_X1 U5921 ( .A(n5865), .B(n5864), .S(n6725), .Z(n5866) );
  MUX2_X1 U5922 ( .A(n5866), .B(n5863), .S(n6709), .Z(n5867) );
  MUX2_X1 U5923 ( .A(n5867), .B(n5860), .S(n6702), .Z(n5868) );
  MUX2_X1 U5924 ( .A(n5868), .B(n5853), .S(addr_r[4]), .Z(n5869) );
  MUX2_X1 U5925 ( .A(n5869), .B(n5838), .S(n6697), .Z(n5870) );
  MUX2_X1 U5926 ( .A(reg_mem[1548]), .B(reg_mem[1540]), .S(n6779), .Z(n5871)
         );
  MUX2_X1 U5927 ( .A(reg_mem[1564]), .B(reg_mem[1556]), .S(n6779), .Z(n5872)
         );
  MUX2_X1 U5928 ( .A(n5872), .B(n5871), .S(n6725), .Z(n5873) );
  MUX2_X1 U5929 ( .A(reg_mem[1580]), .B(reg_mem[1572]), .S(n6779), .Z(n5874)
         );
  MUX2_X1 U5930 ( .A(reg_mem[1596]), .B(reg_mem[1588]), .S(n6770), .Z(n5875)
         );
  MUX2_X1 U5931 ( .A(n5875), .B(n5874), .S(n6725), .Z(n5876) );
  MUX2_X1 U5932 ( .A(n5876), .B(n5873), .S(n6709), .Z(n5877) );
  MUX2_X1 U5933 ( .A(reg_mem[1612]), .B(reg_mem[1604]), .S(n6780), .Z(n5878)
         );
  MUX2_X1 U5934 ( .A(reg_mem[1628]), .B(reg_mem[1620]), .S(n6769), .Z(n5879)
         );
  MUX2_X1 U5935 ( .A(n5879), .B(n5878), .S(n6725), .Z(n5880) );
  MUX2_X1 U5936 ( .A(reg_mem[1644]), .B(reg_mem[1636]), .S(n6771), .Z(n5881)
         );
  MUX2_X1 U5937 ( .A(reg_mem[1660]), .B(reg_mem[1652]), .S(n6773), .Z(n5882)
         );
  MUX2_X1 U5938 ( .A(n5882), .B(n5881), .S(n6725), .Z(n5883) );
  MUX2_X1 U5939 ( .A(n5883), .B(n5880), .S(n6709), .Z(n5884) );
  MUX2_X1 U5940 ( .A(n5884), .B(n5877), .S(n6702), .Z(n5885) );
  MUX2_X1 U5941 ( .A(reg_mem[1676]), .B(reg_mem[1668]), .S(n6749), .Z(n5886)
         );
  MUX2_X1 U5942 ( .A(reg_mem[1692]), .B(reg_mem[1684]), .S(n6749), .Z(n5887)
         );
  MUX2_X1 U5943 ( .A(n5887), .B(n5886), .S(n6719), .Z(n5888) );
  MUX2_X1 U5944 ( .A(reg_mem[1708]), .B(reg_mem[1700]), .S(n6749), .Z(n5889)
         );
  MUX2_X1 U5945 ( .A(reg_mem[1724]), .B(reg_mem[1716]), .S(n6749), .Z(n5890)
         );
  MUX2_X1 U5946 ( .A(n5890), .B(n5889), .S(n6738), .Z(n5891) );
  MUX2_X1 U5947 ( .A(n5891), .B(n5888), .S(n6709), .Z(n5892) );
  MUX2_X1 U5948 ( .A(reg_mem[1740]), .B(reg_mem[1732]), .S(n6749), .Z(n5893)
         );
  MUX2_X1 U5949 ( .A(reg_mem[1756]), .B(reg_mem[1748]), .S(n6749), .Z(n5894)
         );
  MUX2_X1 U5950 ( .A(n5894), .B(n5893), .S(n6737), .Z(n5895) );
  MUX2_X1 U5951 ( .A(reg_mem[1772]), .B(reg_mem[1764]), .S(n6749), .Z(n5896)
         );
  MUX2_X1 U5952 ( .A(reg_mem[1788]), .B(reg_mem[1780]), .S(n6749), .Z(n5897)
         );
  MUX2_X1 U5953 ( .A(n5897), .B(n5896), .S(n6726), .Z(n5898) );
  MUX2_X1 U5954 ( .A(n5898), .B(n5895), .S(n6709), .Z(n5899) );
  MUX2_X1 U5955 ( .A(n5899), .B(n5892), .S(n6702), .Z(n5900) );
  MUX2_X1 U5956 ( .A(n5900), .B(n5885), .S(n6700), .Z(n5901) );
  MUX2_X1 U5957 ( .A(reg_mem[1804]), .B(reg_mem[1796]), .S(n6749), .Z(n5902)
         );
  MUX2_X1 U5958 ( .A(reg_mem[1820]), .B(reg_mem[1812]), .S(n6749), .Z(n5903)
         );
  MUX2_X1 U5959 ( .A(n5903), .B(n5902), .S(n6729), .Z(n5904) );
  MUX2_X1 U5960 ( .A(reg_mem[1836]), .B(reg_mem[1828]), .S(n6749), .Z(n5905)
         );
  MUX2_X1 U5961 ( .A(reg_mem[1852]), .B(reg_mem[1844]), .S(n6749), .Z(n5906)
         );
  MUX2_X1 U5962 ( .A(n5906), .B(n5905), .S(n6730), .Z(n5907) );
  MUX2_X1 U5963 ( .A(n5907), .B(n5904), .S(n6709), .Z(n5908) );
  MUX2_X1 U5964 ( .A(reg_mem[1868]), .B(reg_mem[1860]), .S(n6750), .Z(n5909)
         );
  MUX2_X1 U5965 ( .A(reg_mem[1884]), .B(reg_mem[1876]), .S(n6750), .Z(n5910)
         );
  MUX2_X1 U5966 ( .A(n5910), .B(n5909), .S(n6719), .Z(n5911) );
  MUX2_X1 U5967 ( .A(reg_mem[1900]), .B(reg_mem[1892]), .S(n6750), .Z(n5912)
         );
  MUX2_X1 U5968 ( .A(reg_mem[1916]), .B(reg_mem[1908]), .S(n6750), .Z(n5913)
         );
  MUX2_X1 U5969 ( .A(n5913), .B(n5912), .S(n6727), .Z(n5914) );
  MUX2_X1 U5970 ( .A(n5914), .B(n5911), .S(n6709), .Z(n5915) );
  MUX2_X1 U5971 ( .A(n5915), .B(n5908), .S(n6702), .Z(n5916) );
  MUX2_X1 U5972 ( .A(reg_mem[1932]), .B(reg_mem[1924]), .S(n6750), .Z(n5917)
         );
  MUX2_X1 U5973 ( .A(reg_mem[1948]), .B(reg_mem[1940]), .S(n6750), .Z(n5918)
         );
  MUX2_X1 U5974 ( .A(n5918), .B(n5917), .S(n6738), .Z(n5919) );
  MUX2_X1 U5975 ( .A(reg_mem[1964]), .B(reg_mem[1956]), .S(n6750), .Z(n5920)
         );
  MUX2_X1 U5976 ( .A(reg_mem[1980]), .B(reg_mem[1972]), .S(n6750), .Z(n5921)
         );
  MUX2_X1 U5977 ( .A(n5921), .B(n5920), .S(n6728), .Z(n5922) );
  MUX2_X1 U5978 ( .A(n5922), .B(n5919), .S(n6709), .Z(n5923) );
  MUX2_X1 U5979 ( .A(reg_mem[1996]), .B(reg_mem[1988]), .S(n6750), .Z(n5924)
         );
  MUX2_X1 U5980 ( .A(reg_mem[2012]), .B(reg_mem[2004]), .S(n6750), .Z(n5925)
         );
  MUX2_X1 U5981 ( .A(n5925), .B(n5924), .S(n6738), .Z(n5926) );
  MUX2_X1 U5982 ( .A(reg_mem[2028]), .B(reg_mem[2020]), .S(n6750), .Z(n5927)
         );
  MUX2_X1 U5983 ( .A(reg_mem[2044]), .B(reg_mem[2036]), .S(n6750), .Z(n5928)
         );
  MUX2_X1 U5984 ( .A(n5928), .B(n5927), .S(n6730), .Z(n5929) );
  MUX2_X1 U5985 ( .A(n5929), .B(n5926), .S(n6709), .Z(n5930) );
  MUX2_X1 U5986 ( .A(n5930), .B(n5923), .S(n6702), .Z(n5931) );
  MUX2_X1 U5987 ( .A(n5931), .B(n5916), .S(addr_r[4]), .Z(n5932) );
  MUX2_X1 U5988 ( .A(n5932), .B(n5901), .S(n6697), .Z(n5933) );
  MUX2_X1 U5989 ( .A(n5933), .B(n5870), .S(addr_r[6]), .Z(n5934) );
  MUX2_X1 U5990 ( .A(n5934), .B(n5807), .S(addr_r[7]), .Z(data_r[4]) );
  MUX2_X1 U5991 ( .A(reg_mem[13]), .B(reg_mem[5]), .S(n6751), .Z(n5935) );
  MUX2_X1 U5992 ( .A(reg_mem[29]), .B(reg_mem[21]), .S(n6751), .Z(n5936) );
  MUX2_X1 U5993 ( .A(n5936), .B(n5935), .S(n6730), .Z(n5937) );
  MUX2_X1 U5994 ( .A(reg_mem[45]), .B(reg_mem[37]), .S(n6751), .Z(n5938) );
  MUX2_X1 U5995 ( .A(reg_mem[61]), .B(reg_mem[53]), .S(n6751), .Z(n5939) );
  MUX2_X1 U5996 ( .A(n5939), .B(n5938), .S(n6727), .Z(n5940) );
  MUX2_X1 U5997 ( .A(n5940), .B(n5937), .S(n6710), .Z(n5941) );
  MUX2_X1 U5998 ( .A(reg_mem[77]), .B(reg_mem[69]), .S(n6751), .Z(n5942) );
  MUX2_X1 U5999 ( .A(reg_mem[93]), .B(reg_mem[85]), .S(n6751), .Z(n5943) );
  MUX2_X1 U6000 ( .A(n5943), .B(n5942), .S(n6728), .Z(n5944) );
  MUX2_X1 U6001 ( .A(reg_mem[109]), .B(reg_mem[101]), .S(n6751), .Z(n5945) );
  MUX2_X1 U6002 ( .A(reg_mem[125]), .B(reg_mem[117]), .S(n6751), .Z(n5946) );
  MUX2_X1 U6003 ( .A(n5946), .B(n5945), .S(n6737), .Z(n5947) );
  MUX2_X1 U6004 ( .A(n5947), .B(n5944), .S(n6710), .Z(n5948) );
  MUX2_X1 U6005 ( .A(n5948), .B(n5941), .S(n6703), .Z(n5949) );
  MUX2_X1 U6006 ( .A(reg_mem[141]), .B(reg_mem[133]), .S(n6751), .Z(n5950) );
  MUX2_X1 U6007 ( .A(reg_mem[157]), .B(reg_mem[149]), .S(n6751), .Z(n5951) );
  MUX2_X1 U6008 ( .A(n5951), .B(n5950), .S(n6729), .Z(n5952) );
  MUX2_X1 U6009 ( .A(reg_mem[173]), .B(reg_mem[165]), .S(n6751), .Z(n5953) );
  MUX2_X1 U6010 ( .A(reg_mem[189]), .B(reg_mem[181]), .S(n6751), .Z(n5954) );
  MUX2_X1 U6011 ( .A(n5954), .B(n5953), .S(n6736), .Z(n5955) );
  MUX2_X1 U6012 ( .A(n5955), .B(n5952), .S(n6710), .Z(n5956) );
  MUX2_X1 U6013 ( .A(reg_mem[205]), .B(reg_mem[197]), .S(n6752), .Z(n5957) );
  MUX2_X1 U6014 ( .A(reg_mem[221]), .B(reg_mem[213]), .S(n6752), .Z(n5958) );
  MUX2_X1 U6015 ( .A(n5958), .B(n5957), .S(n6736), .Z(n5959) );
  MUX2_X1 U6016 ( .A(reg_mem[237]), .B(reg_mem[229]), .S(n6752), .Z(n5960) );
  MUX2_X1 U6017 ( .A(reg_mem[253]), .B(reg_mem[245]), .S(n6752), .Z(n5961) );
  MUX2_X1 U6018 ( .A(n5961), .B(n5960), .S(n6728), .Z(n5962) );
  MUX2_X1 U6019 ( .A(n5962), .B(n5959), .S(n6710), .Z(n5963) );
  MUX2_X1 U6020 ( .A(n5963), .B(n5956), .S(n6703), .Z(n5964) );
  MUX2_X1 U6021 ( .A(n5964), .B(n5949), .S(n6698), .Z(n5965) );
  MUX2_X1 U6022 ( .A(reg_mem[269]), .B(reg_mem[261]), .S(n6752), .Z(n5966) );
  MUX2_X1 U6023 ( .A(reg_mem[285]), .B(reg_mem[277]), .S(n6752), .Z(n5967) );
  MUX2_X1 U6024 ( .A(n5967), .B(n5966), .S(n6730), .Z(n5968) );
  MUX2_X1 U6025 ( .A(reg_mem[301]), .B(reg_mem[293]), .S(n6752), .Z(n5969) );
  MUX2_X1 U6026 ( .A(reg_mem[317]), .B(reg_mem[309]), .S(n6752), .Z(n5970) );
  MUX2_X1 U6027 ( .A(n5970), .B(n5969), .S(n6726), .Z(n5971) );
  MUX2_X1 U6028 ( .A(n5971), .B(n5968), .S(n6710), .Z(n5972) );
  MUX2_X1 U6029 ( .A(reg_mem[333]), .B(reg_mem[325]), .S(n6752), .Z(n5973) );
  MUX2_X1 U6030 ( .A(reg_mem[349]), .B(reg_mem[341]), .S(n6752), .Z(n5974) );
  MUX2_X1 U6031 ( .A(n5974), .B(n5973), .S(n6727), .Z(n5975) );
  MUX2_X1 U6032 ( .A(reg_mem[365]), .B(reg_mem[357]), .S(n6752), .Z(n5976) );
  MUX2_X1 U6033 ( .A(reg_mem[381]), .B(reg_mem[373]), .S(n6752), .Z(n5977) );
  MUX2_X1 U6034 ( .A(n5977), .B(n5976), .S(n6729), .Z(n5978) );
  MUX2_X1 U6035 ( .A(n5978), .B(n5975), .S(n6710), .Z(n5979) );
  MUX2_X1 U6036 ( .A(n5979), .B(n5972), .S(n6703), .Z(n5980) );
  MUX2_X1 U6037 ( .A(reg_mem[397]), .B(reg_mem[389]), .S(n6753), .Z(n5981) );
  MUX2_X1 U6038 ( .A(reg_mem[413]), .B(reg_mem[405]), .S(n6753), .Z(n5982) );
  MUX2_X1 U6039 ( .A(n5982), .B(n5981), .S(n6737), .Z(n5983) );
  MUX2_X1 U6040 ( .A(reg_mem[429]), .B(reg_mem[421]), .S(n6753), .Z(n5984) );
  MUX2_X1 U6041 ( .A(reg_mem[445]), .B(reg_mem[437]), .S(n6753), .Z(n5985) );
  MUX2_X1 U6042 ( .A(n5985), .B(n5984), .S(n6737), .Z(n5986) );
  MUX2_X1 U6043 ( .A(n5986), .B(n5983), .S(n6710), .Z(n5987) );
  MUX2_X1 U6044 ( .A(reg_mem[461]), .B(reg_mem[453]), .S(n6753), .Z(n5988) );
  MUX2_X1 U6045 ( .A(reg_mem[477]), .B(reg_mem[469]), .S(n6753), .Z(n5989) );
  MUX2_X1 U6046 ( .A(n5989), .B(n5988), .S(n6738), .Z(n5990) );
  MUX2_X1 U6047 ( .A(reg_mem[493]), .B(reg_mem[485]), .S(n6753), .Z(n5991) );
  MUX2_X1 U6048 ( .A(reg_mem[509]), .B(reg_mem[501]), .S(n6753), .Z(n5992) );
  MUX2_X1 U6049 ( .A(n5992), .B(n5991), .S(n6726), .Z(n5993) );
  MUX2_X1 U6050 ( .A(n5993), .B(n5990), .S(n6710), .Z(n5994) );
  MUX2_X1 U6051 ( .A(n5994), .B(n5987), .S(n6703), .Z(n5995) );
  MUX2_X1 U6052 ( .A(n5995), .B(n5980), .S(n6698), .Z(n5996) );
  MUX2_X1 U6053 ( .A(n5996), .B(n5965), .S(addr_r[5]), .Z(n5997) );
  MUX2_X1 U6054 ( .A(reg_mem[525]), .B(reg_mem[517]), .S(n6753), .Z(n5998) );
  MUX2_X1 U6055 ( .A(reg_mem[541]), .B(reg_mem[533]), .S(n6753), .Z(n5999) );
  MUX2_X1 U6056 ( .A(n5999), .B(n5998), .S(n6725), .Z(n6000) );
  MUX2_X1 U6057 ( .A(reg_mem[557]), .B(reg_mem[549]), .S(n6753), .Z(n6001) );
  MUX2_X1 U6058 ( .A(reg_mem[573]), .B(reg_mem[565]), .S(n6753), .Z(n6002) );
  MUX2_X1 U6059 ( .A(n6002), .B(n6001), .S(n6725), .Z(n6003) );
  MUX2_X1 U6060 ( .A(n6003), .B(n6000), .S(n6710), .Z(n6004) );
  MUX2_X1 U6061 ( .A(reg_mem[589]), .B(reg_mem[581]), .S(n6754), .Z(n6005) );
  MUX2_X1 U6062 ( .A(reg_mem[605]), .B(reg_mem[597]), .S(n6754), .Z(n6006) );
  MUX2_X1 U6063 ( .A(n6006), .B(n6005), .S(n6725), .Z(n6007) );
  MUX2_X1 U6064 ( .A(reg_mem[621]), .B(reg_mem[613]), .S(n6754), .Z(n6008) );
  MUX2_X1 U6065 ( .A(reg_mem[637]), .B(reg_mem[629]), .S(n6754), .Z(n6009) );
  MUX2_X1 U6066 ( .A(n6009), .B(n6008), .S(n6729), .Z(n6010) );
  MUX2_X1 U6067 ( .A(n6010), .B(n6007), .S(n6710), .Z(n6011) );
  MUX2_X1 U6068 ( .A(n6011), .B(n6004), .S(n6703), .Z(n6012) );
  MUX2_X1 U6069 ( .A(reg_mem[653]), .B(reg_mem[645]), .S(n6754), .Z(n6013) );
  MUX2_X1 U6070 ( .A(reg_mem[669]), .B(reg_mem[661]), .S(n6754), .Z(n6014) );
  MUX2_X1 U6071 ( .A(n6014), .B(n6013), .S(n6735), .Z(n6015) );
  MUX2_X1 U6072 ( .A(reg_mem[685]), .B(reg_mem[677]), .S(n6754), .Z(n6016) );
  MUX2_X1 U6073 ( .A(reg_mem[701]), .B(reg_mem[693]), .S(n6754), .Z(n6017) );
  MUX2_X1 U6074 ( .A(n6017), .B(n6016), .S(n6734), .Z(n6018) );
  MUX2_X1 U6075 ( .A(n6018), .B(n6015), .S(n6710), .Z(n6019) );
  MUX2_X1 U6076 ( .A(reg_mem[717]), .B(reg_mem[709]), .S(n6754), .Z(n6020) );
  MUX2_X1 U6077 ( .A(reg_mem[733]), .B(reg_mem[725]), .S(n6754), .Z(n6021) );
  MUX2_X1 U6078 ( .A(n6021), .B(n6020), .S(n6729), .Z(n6022) );
  MUX2_X1 U6079 ( .A(reg_mem[749]), .B(reg_mem[741]), .S(n6754), .Z(n6023) );
  MUX2_X1 U6080 ( .A(reg_mem[765]), .B(reg_mem[757]), .S(n6754), .Z(n6024) );
  MUX2_X1 U6081 ( .A(n6024), .B(n6023), .S(n6726), .Z(n6025) );
  MUX2_X1 U6082 ( .A(n6025), .B(n6022), .S(n6710), .Z(n6026) );
  MUX2_X1 U6083 ( .A(n6026), .B(n6019), .S(n6703), .Z(n6027) );
  MUX2_X1 U6084 ( .A(n6027), .B(n6012), .S(n6698), .Z(n6028) );
  MUX2_X1 U6085 ( .A(reg_mem[781]), .B(reg_mem[773]), .S(n6755), .Z(n6029) );
  MUX2_X1 U6086 ( .A(reg_mem[797]), .B(reg_mem[789]), .S(n6755), .Z(n6030) );
  MUX2_X1 U6087 ( .A(n6030), .B(n6029), .S(n6722), .Z(n6031) );
  MUX2_X1 U6088 ( .A(reg_mem[813]), .B(reg_mem[805]), .S(n6755), .Z(n6032) );
  MUX2_X1 U6089 ( .A(reg_mem[829]), .B(reg_mem[821]), .S(n6755), .Z(n6033) );
  MUX2_X1 U6090 ( .A(n6033), .B(n6032), .S(n6724), .Z(n6034) );
  MUX2_X1 U6091 ( .A(n6034), .B(n6031), .S(n6711), .Z(n6035) );
  MUX2_X1 U6092 ( .A(reg_mem[845]), .B(reg_mem[837]), .S(n6755), .Z(n6036) );
  MUX2_X1 U6093 ( .A(reg_mem[861]), .B(reg_mem[853]), .S(n6755), .Z(n6037) );
  MUX2_X1 U6094 ( .A(n6037), .B(n6036), .S(n6723), .Z(n6038) );
  MUX2_X1 U6095 ( .A(reg_mem[877]), .B(reg_mem[869]), .S(n6755), .Z(n6039) );
  MUX2_X1 U6096 ( .A(reg_mem[893]), .B(reg_mem[885]), .S(n6755), .Z(n6040) );
  MUX2_X1 U6097 ( .A(n6040), .B(n6039), .S(n6738), .Z(n6041) );
  MUX2_X1 U6098 ( .A(n6041), .B(n6038), .S(n6711), .Z(n6042) );
  MUX2_X1 U6099 ( .A(n6042), .B(n6035), .S(n6703), .Z(n6043) );
  MUX2_X1 U6100 ( .A(reg_mem[909]), .B(reg_mem[901]), .S(n6755), .Z(n6044) );
  MUX2_X1 U6101 ( .A(reg_mem[925]), .B(reg_mem[917]), .S(n6755), .Z(n6045) );
  MUX2_X1 U6102 ( .A(n6045), .B(n6044), .S(n6722), .Z(n6046) );
  MUX2_X1 U6103 ( .A(reg_mem[941]), .B(reg_mem[933]), .S(n6755), .Z(n6047) );
  MUX2_X1 U6104 ( .A(reg_mem[957]), .B(reg_mem[949]), .S(n6755), .Z(n6048) );
  MUX2_X1 U6105 ( .A(n6048), .B(n6047), .S(n6724), .Z(n6049) );
  MUX2_X1 U6106 ( .A(n6049), .B(n6046), .S(n6711), .Z(n6050) );
  MUX2_X1 U6107 ( .A(reg_mem[973]), .B(reg_mem[965]), .S(n6756), .Z(n6051) );
  MUX2_X1 U6108 ( .A(reg_mem[989]), .B(reg_mem[981]), .S(n6756), .Z(n6052) );
  MUX2_X1 U6109 ( .A(n6052), .B(n6051), .S(n6723), .Z(n6053) );
  MUX2_X1 U6110 ( .A(reg_mem[1005]), .B(reg_mem[997]), .S(n6756), .Z(n6054) );
  MUX2_X1 U6111 ( .A(reg_mem[1021]), .B(reg_mem[1013]), .S(n6756), .Z(n6055)
         );
  MUX2_X1 U6112 ( .A(n6055), .B(n6054), .S(n6722), .Z(n6056) );
  MUX2_X1 U6113 ( .A(n6056), .B(n6053), .S(n6711), .Z(n6057) );
  MUX2_X1 U6114 ( .A(n6057), .B(n6050), .S(n6703), .Z(n6058) );
  MUX2_X1 U6115 ( .A(n6058), .B(n6043), .S(n6698), .Z(n6059) );
  MUX2_X1 U6116 ( .A(n6059), .B(n6028), .S(n6697), .Z(n6060) );
  MUX2_X1 U6117 ( .A(n6060), .B(n5997), .S(addr_r[6]), .Z(n6061) );
  MUX2_X1 U6118 ( .A(reg_mem[1037]), .B(reg_mem[1029]), .S(n6756), .Z(n6062)
         );
  MUX2_X1 U6119 ( .A(reg_mem[1053]), .B(reg_mem[1045]), .S(n6756), .Z(n6063)
         );
  MUX2_X1 U6120 ( .A(n6063), .B(n6062), .S(n6724), .Z(n6064) );
  MUX2_X1 U6121 ( .A(reg_mem[1069]), .B(reg_mem[1061]), .S(n6756), .Z(n6065)
         );
  MUX2_X1 U6122 ( .A(reg_mem[1085]), .B(reg_mem[1077]), .S(n6756), .Z(n6066)
         );
  MUX2_X1 U6123 ( .A(n6066), .B(n6065), .S(n6724), .Z(n6067) );
  MUX2_X1 U6124 ( .A(n6067), .B(n6064), .S(n6711), .Z(n6068) );
  MUX2_X1 U6125 ( .A(reg_mem[1101]), .B(reg_mem[1093]), .S(n6756), .Z(n6069)
         );
  MUX2_X1 U6126 ( .A(reg_mem[1117]), .B(reg_mem[1109]), .S(n6756), .Z(n6070)
         );
  MUX2_X1 U6127 ( .A(n6070), .B(n6069), .S(n6723), .Z(n6071) );
  MUX2_X1 U6128 ( .A(reg_mem[1133]), .B(reg_mem[1125]), .S(n6756), .Z(n6072)
         );
  MUX2_X1 U6129 ( .A(reg_mem[1149]), .B(reg_mem[1141]), .S(n6756), .Z(n6073)
         );
  MUX2_X1 U6130 ( .A(n6073), .B(n6072), .S(n6730), .Z(n6074) );
  MUX2_X1 U6131 ( .A(n6074), .B(n6071), .S(n6711), .Z(n6075) );
  MUX2_X1 U6132 ( .A(n6075), .B(n6068), .S(n6703), .Z(n6076) );
  MUX2_X1 U6133 ( .A(reg_mem[1165]), .B(reg_mem[1157]), .S(n6757), .Z(n6077)
         );
  MUX2_X1 U6134 ( .A(reg_mem[1181]), .B(reg_mem[1173]), .S(n6757), .Z(n6078)
         );
  MUX2_X1 U6135 ( .A(n6078), .B(n6077), .S(n6726), .Z(n6079) );
  MUX2_X1 U6136 ( .A(reg_mem[1197]), .B(reg_mem[1189]), .S(n6757), .Z(n6080)
         );
  MUX2_X1 U6137 ( .A(reg_mem[1213]), .B(reg_mem[1205]), .S(n6757), .Z(n6081)
         );
  MUX2_X1 U6138 ( .A(n6081), .B(n6080), .S(n6726), .Z(n6082) );
  MUX2_X1 U6139 ( .A(n6082), .B(n6079), .S(n6711), .Z(n6083) );
  MUX2_X1 U6140 ( .A(reg_mem[1229]), .B(reg_mem[1221]), .S(n6757), .Z(n6084)
         );
  MUX2_X1 U6141 ( .A(reg_mem[1245]), .B(reg_mem[1237]), .S(n6757), .Z(n6085)
         );
  MUX2_X1 U6142 ( .A(n6085), .B(n6084), .S(n6726), .Z(n6086) );
  MUX2_X1 U6143 ( .A(reg_mem[1261]), .B(reg_mem[1253]), .S(n6757), .Z(n6087)
         );
  MUX2_X1 U6144 ( .A(reg_mem[1277]), .B(reg_mem[1269]), .S(n6757), .Z(n6088)
         );
  MUX2_X1 U6145 ( .A(n6088), .B(n6087), .S(n6726), .Z(n6089) );
  MUX2_X1 U6146 ( .A(n6089), .B(n6086), .S(n6711), .Z(n6090) );
  MUX2_X1 U6147 ( .A(n6090), .B(n6083), .S(n6703), .Z(n6091) );
  MUX2_X1 U6148 ( .A(n6091), .B(n6076), .S(n6698), .Z(n6092) );
  MUX2_X1 U6149 ( .A(reg_mem[1293]), .B(reg_mem[1285]), .S(n6757), .Z(n6093)
         );
  MUX2_X1 U6150 ( .A(reg_mem[1309]), .B(reg_mem[1301]), .S(n6757), .Z(n6094)
         );
  MUX2_X1 U6151 ( .A(n6094), .B(n6093), .S(n6726), .Z(n6095) );
  MUX2_X1 U6152 ( .A(reg_mem[1325]), .B(reg_mem[1317]), .S(n6757), .Z(n6096)
         );
  MUX2_X1 U6153 ( .A(reg_mem[1341]), .B(reg_mem[1333]), .S(n6757), .Z(n6097)
         );
  MUX2_X1 U6154 ( .A(n6097), .B(n6096), .S(n6726), .Z(n6098) );
  MUX2_X1 U6155 ( .A(n6098), .B(n6095), .S(n6711), .Z(n6099) );
  MUX2_X1 U6156 ( .A(reg_mem[1357]), .B(reg_mem[1349]), .S(n6758), .Z(n6100)
         );
  MUX2_X1 U6157 ( .A(reg_mem[1373]), .B(reg_mem[1365]), .S(n6758), .Z(n6101)
         );
  MUX2_X1 U6158 ( .A(n6101), .B(n6100), .S(n6726), .Z(n6102) );
  MUX2_X1 U6159 ( .A(reg_mem[1389]), .B(reg_mem[1381]), .S(n6758), .Z(n6103)
         );
  MUX2_X1 U6160 ( .A(reg_mem[1405]), .B(reg_mem[1397]), .S(n6758), .Z(n6104)
         );
  MUX2_X1 U6161 ( .A(n6104), .B(n6103), .S(n6726), .Z(n6105) );
  MUX2_X1 U6162 ( .A(n6105), .B(n6102), .S(n6711), .Z(n6106) );
  MUX2_X1 U6163 ( .A(n6106), .B(n6099), .S(n6703), .Z(n6107) );
  MUX2_X1 U6164 ( .A(reg_mem[1421]), .B(reg_mem[1413]), .S(n6758), .Z(n6108)
         );
  MUX2_X1 U6165 ( .A(reg_mem[1437]), .B(reg_mem[1429]), .S(n6758), .Z(n6109)
         );
  MUX2_X1 U6166 ( .A(n6109), .B(n6108), .S(n6726), .Z(n6110) );
  MUX2_X1 U6167 ( .A(reg_mem[1453]), .B(reg_mem[1445]), .S(n6758), .Z(n6111)
         );
  MUX2_X1 U6168 ( .A(reg_mem[1469]), .B(reg_mem[1461]), .S(n6758), .Z(n6112)
         );
  MUX2_X1 U6169 ( .A(n6112), .B(n6111), .S(n6726), .Z(n6113) );
  MUX2_X1 U6170 ( .A(n6113), .B(n6110), .S(n6711), .Z(n6114) );
  MUX2_X1 U6171 ( .A(reg_mem[1485]), .B(reg_mem[1477]), .S(n6758), .Z(n6115)
         );
  MUX2_X1 U6172 ( .A(reg_mem[1501]), .B(reg_mem[1493]), .S(n6758), .Z(n6116)
         );
  MUX2_X1 U6173 ( .A(n6116), .B(n6115), .S(n6726), .Z(n6117) );
  MUX2_X1 U6174 ( .A(reg_mem[1517]), .B(reg_mem[1509]), .S(n6758), .Z(n6118)
         );
  MUX2_X1 U6175 ( .A(reg_mem[1533]), .B(reg_mem[1525]), .S(n6758), .Z(n6119)
         );
  MUX2_X1 U6176 ( .A(n6119), .B(n6118), .S(n6726), .Z(n6120) );
  MUX2_X1 U6177 ( .A(n6120), .B(n6117), .S(n6711), .Z(n6121) );
  MUX2_X1 U6178 ( .A(n6121), .B(n6114), .S(n6703), .Z(n6122) );
  MUX2_X1 U6179 ( .A(n6122), .B(n6107), .S(n6698), .Z(n6123) );
  MUX2_X1 U6180 ( .A(n6123), .B(n6092), .S(n6697), .Z(n6124) );
  MUX2_X1 U6181 ( .A(reg_mem[1549]), .B(reg_mem[1541]), .S(n6759), .Z(n6125)
         );
  MUX2_X1 U6182 ( .A(reg_mem[1565]), .B(reg_mem[1557]), .S(n6759), .Z(n6126)
         );
  MUX2_X1 U6183 ( .A(n6126), .B(n6125), .S(n6727), .Z(n6127) );
  MUX2_X1 U6184 ( .A(reg_mem[1581]), .B(reg_mem[1573]), .S(n6759), .Z(n6128)
         );
  MUX2_X1 U6185 ( .A(reg_mem[1597]), .B(reg_mem[1589]), .S(n6759), .Z(n6129)
         );
  MUX2_X1 U6186 ( .A(n6129), .B(n6128), .S(n6727), .Z(n6130) );
  MUX2_X1 U6187 ( .A(n6130), .B(n6127), .S(n6712), .Z(n6131) );
  MUX2_X1 U6188 ( .A(reg_mem[1613]), .B(reg_mem[1605]), .S(n6759), .Z(n6132)
         );
  MUX2_X1 U6189 ( .A(reg_mem[1629]), .B(reg_mem[1621]), .S(n6759), .Z(n6133)
         );
  MUX2_X1 U6190 ( .A(n6133), .B(n6132), .S(n6727), .Z(n6134) );
  MUX2_X1 U6191 ( .A(reg_mem[1645]), .B(reg_mem[1637]), .S(n6759), .Z(n6135)
         );
  MUX2_X1 U6192 ( .A(reg_mem[1661]), .B(reg_mem[1653]), .S(n6759), .Z(n6136)
         );
  MUX2_X1 U6193 ( .A(n6136), .B(n6135), .S(n6727), .Z(n6137) );
  MUX2_X1 U6194 ( .A(n6137), .B(n6134), .S(n6712), .Z(n6138) );
  MUX2_X1 U6195 ( .A(n6138), .B(n6131), .S(n6704), .Z(n6139) );
  MUX2_X1 U6196 ( .A(reg_mem[1677]), .B(reg_mem[1669]), .S(n6759), .Z(n6140)
         );
  MUX2_X1 U6197 ( .A(reg_mem[1693]), .B(reg_mem[1685]), .S(n6759), .Z(n6141)
         );
  MUX2_X1 U6198 ( .A(n6141), .B(n6140), .S(n6727), .Z(n6142) );
  MUX2_X1 U6199 ( .A(reg_mem[1709]), .B(reg_mem[1701]), .S(n6759), .Z(n6143)
         );
  MUX2_X1 U6200 ( .A(reg_mem[1725]), .B(reg_mem[1717]), .S(n6759), .Z(n6144)
         );
  MUX2_X1 U6201 ( .A(n6144), .B(n6143), .S(n6727), .Z(n6145) );
  MUX2_X1 U6202 ( .A(n6145), .B(n6142), .S(n6712), .Z(n6146) );
  MUX2_X1 U6203 ( .A(reg_mem[1741]), .B(reg_mem[1733]), .S(n6760), .Z(n6147)
         );
  MUX2_X1 U6204 ( .A(reg_mem[1757]), .B(reg_mem[1749]), .S(n6760), .Z(n6148)
         );
  MUX2_X1 U6205 ( .A(n6148), .B(n6147), .S(n6727), .Z(n6149) );
  MUX2_X1 U6206 ( .A(reg_mem[1773]), .B(reg_mem[1765]), .S(n6760), .Z(n6150)
         );
  MUX2_X1 U6207 ( .A(reg_mem[1789]), .B(reg_mem[1781]), .S(n6760), .Z(n6151)
         );
  MUX2_X1 U6208 ( .A(n6151), .B(n6150), .S(n6727), .Z(n6152) );
  MUX2_X1 U6209 ( .A(n6152), .B(n6149), .S(n6712), .Z(n6153) );
  MUX2_X1 U6210 ( .A(n6153), .B(n6146), .S(n6704), .Z(n6154) );
  MUX2_X1 U6211 ( .A(n6154), .B(n6139), .S(n6698), .Z(n6155) );
  MUX2_X1 U6212 ( .A(reg_mem[1805]), .B(reg_mem[1797]), .S(n6760), .Z(n6156)
         );
  MUX2_X1 U6213 ( .A(reg_mem[1821]), .B(reg_mem[1813]), .S(n6760), .Z(n6157)
         );
  MUX2_X1 U6214 ( .A(n6157), .B(n6156), .S(n6727), .Z(n6158) );
  MUX2_X1 U6215 ( .A(reg_mem[1837]), .B(reg_mem[1829]), .S(n6760), .Z(n6159)
         );
  MUX2_X1 U6216 ( .A(reg_mem[1853]), .B(reg_mem[1845]), .S(n6760), .Z(n6160)
         );
  MUX2_X1 U6217 ( .A(n6160), .B(n6159), .S(n6727), .Z(n6161) );
  MUX2_X1 U6218 ( .A(n6161), .B(n6158), .S(n6712), .Z(n6162) );
  MUX2_X1 U6219 ( .A(reg_mem[1869]), .B(reg_mem[1861]), .S(n6760), .Z(n6163)
         );
  MUX2_X1 U6220 ( .A(reg_mem[1885]), .B(reg_mem[1877]), .S(n6760), .Z(n6164)
         );
  MUX2_X1 U6221 ( .A(n6164), .B(n6163), .S(n6727), .Z(n6165) );
  MUX2_X1 U6222 ( .A(reg_mem[1901]), .B(reg_mem[1893]), .S(n6760), .Z(n6166)
         );
  MUX2_X1 U6223 ( .A(reg_mem[1917]), .B(reg_mem[1909]), .S(n6760), .Z(n6167)
         );
  MUX2_X1 U6224 ( .A(n6167), .B(n6166), .S(n6727), .Z(n6168) );
  MUX2_X1 U6225 ( .A(n6168), .B(n6165), .S(n6712), .Z(n6169) );
  MUX2_X1 U6226 ( .A(n6169), .B(n6162), .S(n6704), .Z(n6170) );
  MUX2_X1 U6227 ( .A(reg_mem[1933]), .B(reg_mem[1925]), .S(n6761), .Z(n6171)
         );
  MUX2_X1 U6228 ( .A(reg_mem[1949]), .B(reg_mem[1941]), .S(n6761), .Z(n6172)
         );
  MUX2_X1 U6229 ( .A(n6172), .B(n6171), .S(n6728), .Z(n6173) );
  MUX2_X1 U6230 ( .A(reg_mem[1965]), .B(reg_mem[1957]), .S(n6761), .Z(n6174)
         );
  MUX2_X1 U6231 ( .A(reg_mem[1981]), .B(reg_mem[1973]), .S(n6761), .Z(n6175)
         );
  MUX2_X1 U6232 ( .A(n6175), .B(n6174), .S(n6728), .Z(n6176) );
  MUX2_X1 U6233 ( .A(n6176), .B(n6173), .S(n6712), .Z(n6177) );
  MUX2_X1 U6234 ( .A(reg_mem[1997]), .B(reg_mem[1989]), .S(n6761), .Z(n6178)
         );
  MUX2_X1 U6235 ( .A(reg_mem[2013]), .B(reg_mem[2005]), .S(n6761), .Z(n6179)
         );
  MUX2_X1 U6236 ( .A(n6179), .B(n6178), .S(n6728), .Z(n6180) );
  MUX2_X1 U6237 ( .A(reg_mem[2029]), .B(reg_mem[2021]), .S(n6761), .Z(n6181)
         );
  MUX2_X1 U6238 ( .A(reg_mem[2045]), .B(reg_mem[2037]), .S(n6761), .Z(n6182)
         );
  MUX2_X1 U6239 ( .A(n6182), .B(n6181), .S(n6728), .Z(n6183) );
  MUX2_X1 U6240 ( .A(n6183), .B(n6180), .S(n6712), .Z(n6184) );
  MUX2_X1 U6241 ( .A(n6184), .B(n6177), .S(n6704), .Z(n6185) );
  MUX2_X1 U6242 ( .A(n6185), .B(n6170), .S(n6698), .Z(n6186) );
  MUX2_X1 U6243 ( .A(n6186), .B(n6155), .S(n6697), .Z(n6187) );
  MUX2_X1 U6244 ( .A(n6187), .B(n6124), .S(addr_r[6]), .Z(n6188) );
  MUX2_X1 U6245 ( .A(n6188), .B(n6061), .S(addr_r[7]), .Z(data_r[5]) );
  MUX2_X1 U6246 ( .A(reg_mem[14]), .B(reg_mem[6]), .S(n6761), .Z(n6189) );
  MUX2_X1 U6247 ( .A(reg_mem[30]), .B(reg_mem[22]), .S(n6761), .Z(n6190) );
  MUX2_X1 U6248 ( .A(n6190), .B(n6189), .S(n6728), .Z(n6191) );
  MUX2_X1 U6249 ( .A(reg_mem[46]), .B(reg_mem[38]), .S(n6761), .Z(n6192) );
  MUX2_X1 U6250 ( .A(reg_mem[62]), .B(reg_mem[54]), .S(n6761), .Z(n6193) );
  MUX2_X1 U6251 ( .A(n6193), .B(n6192), .S(n6728), .Z(n6194) );
  MUX2_X1 U6252 ( .A(n6194), .B(n6191), .S(n6712), .Z(n6195) );
  MUX2_X1 U6253 ( .A(reg_mem[78]), .B(reg_mem[70]), .S(n6762), .Z(n6196) );
  MUX2_X1 U6254 ( .A(reg_mem[94]), .B(reg_mem[86]), .S(n6762), .Z(n6197) );
  MUX2_X1 U6255 ( .A(n6197), .B(n6196), .S(n6728), .Z(n6198) );
  MUX2_X1 U6256 ( .A(reg_mem[110]), .B(reg_mem[102]), .S(n6762), .Z(n6199) );
  MUX2_X1 U6257 ( .A(reg_mem[126]), .B(reg_mem[118]), .S(n6762), .Z(n6200) );
  MUX2_X1 U6258 ( .A(n6200), .B(n6199), .S(n6728), .Z(n6201) );
  MUX2_X1 U6259 ( .A(n6201), .B(n6198), .S(n6712), .Z(n6202) );
  MUX2_X1 U6260 ( .A(n6202), .B(n6195), .S(n6704), .Z(n6203) );
  MUX2_X1 U6261 ( .A(reg_mem[142]), .B(reg_mem[134]), .S(n6762), .Z(n6204) );
  MUX2_X1 U6262 ( .A(reg_mem[158]), .B(reg_mem[150]), .S(n6762), .Z(n6205) );
  MUX2_X1 U6263 ( .A(n6205), .B(n6204), .S(n6728), .Z(n6206) );
  MUX2_X1 U6264 ( .A(reg_mem[174]), .B(reg_mem[166]), .S(n6762), .Z(n6207) );
  MUX2_X1 U6265 ( .A(reg_mem[190]), .B(reg_mem[182]), .S(n6762), .Z(n6208) );
  MUX2_X1 U6266 ( .A(n6208), .B(n6207), .S(n6728), .Z(n6209) );
  MUX2_X1 U6267 ( .A(n6209), .B(n6206), .S(n6712), .Z(n6210) );
  MUX2_X1 U6268 ( .A(reg_mem[206]), .B(reg_mem[198]), .S(n6762), .Z(n6211) );
  MUX2_X1 U6269 ( .A(reg_mem[222]), .B(reg_mem[214]), .S(n6762), .Z(n6212) );
  MUX2_X1 U6270 ( .A(n6212), .B(n6211), .S(n6728), .Z(n6213) );
  MUX2_X1 U6271 ( .A(reg_mem[238]), .B(reg_mem[230]), .S(n6762), .Z(n6214) );
  MUX2_X1 U6272 ( .A(reg_mem[254]), .B(reg_mem[246]), .S(n6762), .Z(n6215) );
  MUX2_X1 U6273 ( .A(n6215), .B(n6214), .S(n6728), .Z(n6216) );
  MUX2_X1 U6274 ( .A(n6216), .B(n6213), .S(n6712), .Z(n6217) );
  MUX2_X1 U6275 ( .A(n6217), .B(n6210), .S(n6704), .Z(n6218) );
  MUX2_X1 U6276 ( .A(n6218), .B(n6203), .S(n6698), .Z(n6219) );
  MUX2_X1 U6277 ( .A(reg_mem[270]), .B(reg_mem[262]), .S(n6763), .Z(n6220) );
  MUX2_X1 U6278 ( .A(reg_mem[286]), .B(reg_mem[278]), .S(n6763), .Z(n6221) );
  MUX2_X1 U6279 ( .A(n6221), .B(n6220), .S(n6729), .Z(n6222) );
  MUX2_X1 U6280 ( .A(reg_mem[302]), .B(reg_mem[294]), .S(n6763), .Z(n6223) );
  MUX2_X1 U6281 ( .A(reg_mem[318]), .B(reg_mem[310]), .S(n6763), .Z(n6224) );
  MUX2_X1 U6282 ( .A(n6224), .B(n6223), .S(n6729), .Z(n6225) );
  MUX2_X1 U6283 ( .A(n6225), .B(n6222), .S(n6713), .Z(n6226) );
  MUX2_X1 U6284 ( .A(reg_mem[334]), .B(reg_mem[326]), .S(n6763), .Z(n6227) );
  MUX2_X1 U6285 ( .A(reg_mem[350]), .B(reg_mem[342]), .S(n6763), .Z(n6228) );
  MUX2_X1 U6286 ( .A(n6228), .B(n6227), .S(n6729), .Z(n6229) );
  MUX2_X1 U6287 ( .A(reg_mem[366]), .B(reg_mem[358]), .S(n6763), .Z(n6230) );
  MUX2_X1 U6288 ( .A(reg_mem[382]), .B(reg_mem[374]), .S(n6763), .Z(n6231) );
  MUX2_X1 U6289 ( .A(n6231), .B(n6230), .S(n6729), .Z(n6232) );
  MUX2_X1 U6290 ( .A(n6232), .B(n6229), .S(n6713), .Z(n6233) );
  MUX2_X1 U6291 ( .A(n6233), .B(n6226), .S(n6704), .Z(n6234) );
  MUX2_X1 U6292 ( .A(reg_mem[398]), .B(reg_mem[390]), .S(n6763), .Z(n6235) );
  MUX2_X1 U6293 ( .A(reg_mem[414]), .B(reg_mem[406]), .S(n6763), .Z(n6236) );
  MUX2_X1 U6294 ( .A(n6236), .B(n6235), .S(n6729), .Z(n6237) );
  MUX2_X1 U6295 ( .A(reg_mem[430]), .B(reg_mem[422]), .S(n6763), .Z(n6238) );
  MUX2_X1 U6296 ( .A(reg_mem[446]), .B(reg_mem[438]), .S(n6763), .Z(n6239) );
  MUX2_X1 U6297 ( .A(n6239), .B(n6238), .S(n6729), .Z(n6240) );
  MUX2_X1 U6298 ( .A(n6240), .B(n6237), .S(n6713), .Z(n6241) );
  MUX2_X1 U6299 ( .A(reg_mem[462]), .B(reg_mem[454]), .S(n6764), .Z(n6242) );
  MUX2_X1 U6300 ( .A(reg_mem[478]), .B(reg_mem[470]), .S(n6764), .Z(n6243) );
  MUX2_X1 U6301 ( .A(n6243), .B(n6242), .S(n6729), .Z(n6244) );
  MUX2_X1 U6302 ( .A(reg_mem[494]), .B(reg_mem[486]), .S(n6764), .Z(n6245) );
  MUX2_X1 U6303 ( .A(reg_mem[510]), .B(reg_mem[502]), .S(n6764), .Z(n6246) );
  MUX2_X1 U6304 ( .A(n6246), .B(n6245), .S(n6729), .Z(n6247) );
  MUX2_X1 U6305 ( .A(n6247), .B(n6244), .S(n6713), .Z(n6248) );
  MUX2_X1 U6306 ( .A(n6248), .B(n6241), .S(n6704), .Z(n6249) );
  MUX2_X1 U6307 ( .A(n6249), .B(n6234), .S(n6698), .Z(n6250) );
  MUX2_X1 U6308 ( .A(n6250), .B(n6219), .S(addr_r[5]), .Z(n6251) );
  MUX2_X1 U6309 ( .A(reg_mem[526]), .B(reg_mem[518]), .S(n6764), .Z(n6252) );
  MUX2_X1 U6310 ( .A(reg_mem[542]), .B(reg_mem[534]), .S(n6764), .Z(n6253) );
  MUX2_X1 U6311 ( .A(n6253), .B(n6252), .S(n6729), .Z(n6254) );
  MUX2_X1 U6312 ( .A(reg_mem[558]), .B(reg_mem[550]), .S(n6764), .Z(n6255) );
  MUX2_X1 U6313 ( .A(reg_mem[574]), .B(reg_mem[566]), .S(n6764), .Z(n6256) );
  MUX2_X1 U6314 ( .A(n6256), .B(n6255), .S(n6729), .Z(n6257) );
  MUX2_X1 U6315 ( .A(n6257), .B(n6254), .S(n6713), .Z(n6258) );
  MUX2_X1 U6316 ( .A(reg_mem[590]), .B(reg_mem[582]), .S(n6764), .Z(n6259) );
  MUX2_X1 U6317 ( .A(reg_mem[606]), .B(reg_mem[598]), .S(n6764), .Z(n6260) );
  MUX2_X1 U6318 ( .A(n6260), .B(n6259), .S(n6729), .Z(n6261) );
  MUX2_X1 U6319 ( .A(reg_mem[622]), .B(reg_mem[614]), .S(n6764), .Z(n6262) );
  MUX2_X1 U6320 ( .A(reg_mem[638]), .B(reg_mem[630]), .S(n6764), .Z(n6263) );
  MUX2_X1 U6321 ( .A(n6263), .B(n6262), .S(n6729), .Z(n6264) );
  MUX2_X1 U6322 ( .A(n6264), .B(n6261), .S(n6713), .Z(n6265) );
  MUX2_X1 U6323 ( .A(n6265), .B(n6258), .S(n6704), .Z(n6266) );
  MUX2_X1 U6324 ( .A(reg_mem[654]), .B(reg_mem[646]), .S(n6765), .Z(n6267) );
  MUX2_X1 U6325 ( .A(reg_mem[670]), .B(reg_mem[662]), .S(n6765), .Z(n6268) );
  MUX2_X1 U6326 ( .A(n6268), .B(n6267), .S(n6730), .Z(n6269) );
  MUX2_X1 U6327 ( .A(reg_mem[686]), .B(reg_mem[678]), .S(n6765), .Z(n6270) );
  MUX2_X1 U6328 ( .A(reg_mem[702]), .B(reg_mem[694]), .S(n6765), .Z(n6271) );
  MUX2_X1 U6329 ( .A(n6271), .B(n6270), .S(n6730), .Z(n6272) );
  MUX2_X1 U6330 ( .A(n6272), .B(n6269), .S(n6713), .Z(n6273) );
  MUX2_X1 U6331 ( .A(reg_mem[718]), .B(reg_mem[710]), .S(n6765), .Z(n6274) );
  MUX2_X1 U6332 ( .A(reg_mem[734]), .B(reg_mem[726]), .S(n6765), .Z(n6275) );
  MUX2_X1 U6333 ( .A(n6275), .B(n6274), .S(n6730), .Z(n6276) );
  MUX2_X1 U6334 ( .A(reg_mem[750]), .B(reg_mem[742]), .S(n6765), .Z(n6277) );
  MUX2_X1 U6335 ( .A(reg_mem[766]), .B(reg_mem[758]), .S(n6765), .Z(n6278) );
  MUX2_X1 U6336 ( .A(n6278), .B(n6277), .S(n6730), .Z(n6279) );
  MUX2_X1 U6337 ( .A(n6279), .B(n6276), .S(n6713), .Z(n6280) );
  MUX2_X1 U6338 ( .A(n6280), .B(n6273), .S(n6704), .Z(n6281) );
  MUX2_X1 U6339 ( .A(n6281), .B(n6266), .S(n6698), .Z(n6282) );
  MUX2_X1 U6340 ( .A(reg_mem[782]), .B(reg_mem[774]), .S(n6765), .Z(n6283) );
  MUX2_X1 U6341 ( .A(reg_mem[798]), .B(reg_mem[790]), .S(n6765), .Z(n6284) );
  MUX2_X1 U6342 ( .A(n6284), .B(n6283), .S(n6730), .Z(n6285) );
  MUX2_X1 U6343 ( .A(reg_mem[814]), .B(reg_mem[806]), .S(n6765), .Z(n6286) );
  MUX2_X1 U6344 ( .A(reg_mem[830]), .B(reg_mem[822]), .S(n6765), .Z(n6287) );
  MUX2_X1 U6345 ( .A(n6287), .B(n6286), .S(n6730), .Z(n6288) );
  MUX2_X1 U6346 ( .A(n6288), .B(n6285), .S(n6713), .Z(n6289) );
  MUX2_X1 U6347 ( .A(reg_mem[846]), .B(reg_mem[838]), .S(n6766), .Z(n6290) );
  MUX2_X1 U6348 ( .A(reg_mem[862]), .B(reg_mem[854]), .S(n6766), .Z(n6291) );
  MUX2_X1 U6349 ( .A(n6291), .B(n6290), .S(n6730), .Z(n6292) );
  MUX2_X1 U6350 ( .A(reg_mem[878]), .B(reg_mem[870]), .S(n6766), .Z(n6293) );
  MUX2_X1 U6351 ( .A(reg_mem[894]), .B(reg_mem[886]), .S(n6766), .Z(n6294) );
  MUX2_X1 U6352 ( .A(n6294), .B(n6293), .S(n6730), .Z(n6295) );
  MUX2_X1 U6353 ( .A(n6295), .B(n6292), .S(n6713), .Z(n6296) );
  MUX2_X1 U6354 ( .A(n6296), .B(n6289), .S(n6704), .Z(n6297) );
  MUX2_X1 U6355 ( .A(reg_mem[910]), .B(reg_mem[902]), .S(n6766), .Z(n6298) );
  MUX2_X1 U6356 ( .A(reg_mem[926]), .B(reg_mem[918]), .S(n6766), .Z(n6299) );
  MUX2_X1 U6357 ( .A(n6299), .B(n6298), .S(n6730), .Z(n6300) );
  MUX2_X1 U6358 ( .A(reg_mem[942]), .B(reg_mem[934]), .S(n6766), .Z(n6301) );
  MUX2_X1 U6359 ( .A(reg_mem[958]), .B(reg_mem[950]), .S(n6766), .Z(n6302) );
  MUX2_X1 U6360 ( .A(n6302), .B(n6301), .S(n6730), .Z(n6303) );
  MUX2_X1 U6361 ( .A(n6303), .B(n6300), .S(n6713), .Z(n6304) );
  MUX2_X1 U6362 ( .A(reg_mem[974]), .B(reg_mem[966]), .S(n6766), .Z(n6305) );
  MUX2_X1 U6363 ( .A(reg_mem[990]), .B(reg_mem[982]), .S(n6766), .Z(n6306) );
  MUX2_X1 U6364 ( .A(n6306), .B(n6305), .S(n6730), .Z(n6307) );
  MUX2_X1 U6365 ( .A(reg_mem[1006]), .B(reg_mem[998]), .S(n6766), .Z(n6308) );
  MUX2_X1 U6366 ( .A(reg_mem[1022]), .B(reg_mem[1014]), .S(n6766), .Z(n6309)
         );
  MUX2_X1 U6367 ( .A(n6309), .B(n6308), .S(n6730), .Z(n6310) );
  MUX2_X1 U6368 ( .A(n6310), .B(n6307), .S(n6713), .Z(n6311) );
  MUX2_X1 U6369 ( .A(n6311), .B(n6304), .S(n6704), .Z(n6312) );
  MUX2_X1 U6370 ( .A(n6312), .B(n6297), .S(n6698), .Z(n6313) );
  MUX2_X1 U6371 ( .A(n6313), .B(n6282), .S(n6697), .Z(n6314) );
  MUX2_X1 U6372 ( .A(n6314), .B(n6251), .S(addr_r[6]), .Z(n6315) );
  MUX2_X1 U6373 ( .A(reg_mem[1038]), .B(reg_mem[1030]), .S(n6767), .Z(n6316)
         );
  MUX2_X1 U6374 ( .A(reg_mem[1054]), .B(reg_mem[1046]), .S(n6767), .Z(n6317)
         );
  MUX2_X1 U6375 ( .A(n6317), .B(n6316), .S(n6731), .Z(n6318) );
  MUX2_X1 U6376 ( .A(reg_mem[1070]), .B(reg_mem[1062]), .S(n6767), .Z(n6319)
         );
  MUX2_X1 U6377 ( .A(reg_mem[1086]), .B(reg_mem[1078]), .S(n6767), .Z(n6320)
         );
  MUX2_X1 U6378 ( .A(n6320), .B(n6319), .S(n6731), .Z(n6321) );
  MUX2_X1 U6379 ( .A(n6321), .B(n6318), .S(n6714), .Z(n6322) );
  MUX2_X1 U6380 ( .A(reg_mem[1102]), .B(reg_mem[1094]), .S(n6767), .Z(n6323)
         );
  MUX2_X1 U6381 ( .A(reg_mem[1118]), .B(reg_mem[1110]), .S(n6767), .Z(n6324)
         );
  MUX2_X1 U6382 ( .A(n6324), .B(n6323), .S(n6731), .Z(n6325) );
  MUX2_X1 U6383 ( .A(reg_mem[1134]), .B(reg_mem[1126]), .S(n6767), .Z(n6326)
         );
  MUX2_X1 U6384 ( .A(reg_mem[1150]), .B(reg_mem[1142]), .S(n6767), .Z(n6327)
         );
  MUX2_X1 U6385 ( .A(n6327), .B(n6326), .S(n6731), .Z(n6328) );
  MUX2_X1 U6386 ( .A(n6328), .B(n6325), .S(n6714), .Z(n6329) );
  MUX2_X1 U6387 ( .A(n6329), .B(n6322), .S(n6705), .Z(n6330) );
  MUX2_X1 U6388 ( .A(reg_mem[1166]), .B(reg_mem[1158]), .S(n6767), .Z(n6331)
         );
  MUX2_X1 U6389 ( .A(reg_mem[1182]), .B(reg_mem[1174]), .S(n6767), .Z(n6332)
         );
  MUX2_X1 U6390 ( .A(n6332), .B(n6331), .S(n6731), .Z(n6333) );
  MUX2_X1 U6391 ( .A(reg_mem[1198]), .B(reg_mem[1190]), .S(n6767), .Z(n6334)
         );
  MUX2_X1 U6392 ( .A(reg_mem[1214]), .B(reg_mem[1206]), .S(n6767), .Z(n6335)
         );
  MUX2_X1 U6393 ( .A(n6335), .B(n6334), .S(n6731), .Z(n6336) );
  MUX2_X1 U6394 ( .A(n6336), .B(n6333), .S(n6714), .Z(n6337) );
  MUX2_X1 U6395 ( .A(reg_mem[1230]), .B(reg_mem[1222]), .S(n6768), .Z(n6338)
         );
  MUX2_X1 U6396 ( .A(reg_mem[1246]), .B(reg_mem[1238]), .S(n6768), .Z(n6339)
         );
  MUX2_X1 U6397 ( .A(n6339), .B(n6338), .S(n6731), .Z(n6340) );
  MUX2_X1 U6398 ( .A(reg_mem[1262]), .B(reg_mem[1254]), .S(n6768), .Z(n6341)
         );
  MUX2_X1 U6399 ( .A(reg_mem[1278]), .B(reg_mem[1270]), .S(n6768), .Z(n6342)
         );
  MUX2_X1 U6400 ( .A(n6342), .B(n6341), .S(n6731), .Z(n6343) );
  MUX2_X1 U6401 ( .A(n6343), .B(n6340), .S(n6714), .Z(n6344) );
  MUX2_X1 U6402 ( .A(n6344), .B(n6337), .S(n6705), .Z(n6345) );
  MUX2_X1 U6403 ( .A(n6345), .B(n6330), .S(n6699), .Z(n6346) );
  MUX2_X1 U6404 ( .A(reg_mem[1294]), .B(reg_mem[1286]), .S(n6768), .Z(n6347)
         );
  MUX2_X1 U6405 ( .A(reg_mem[1310]), .B(reg_mem[1302]), .S(n6768), .Z(n6348)
         );
  MUX2_X1 U6406 ( .A(n6348), .B(n6347), .S(n6731), .Z(n6349) );
  MUX2_X1 U6407 ( .A(reg_mem[1326]), .B(reg_mem[1318]), .S(n6768), .Z(n6350)
         );
  MUX2_X1 U6408 ( .A(reg_mem[1342]), .B(reg_mem[1334]), .S(n6768), .Z(n6351)
         );
  MUX2_X1 U6409 ( .A(n6351), .B(n6350), .S(n6731), .Z(n6352) );
  MUX2_X1 U6410 ( .A(n6352), .B(n6349), .S(n6714), .Z(n6353) );
  MUX2_X1 U6411 ( .A(reg_mem[1358]), .B(reg_mem[1350]), .S(n6768), .Z(n6354)
         );
  MUX2_X1 U6412 ( .A(reg_mem[1374]), .B(reg_mem[1366]), .S(n6768), .Z(n6355)
         );
  MUX2_X1 U6413 ( .A(n6355), .B(n6354), .S(n6731), .Z(n6356) );
  MUX2_X1 U6414 ( .A(reg_mem[1390]), .B(reg_mem[1382]), .S(n6768), .Z(n6357)
         );
  MUX2_X1 U6415 ( .A(reg_mem[1406]), .B(reg_mem[1398]), .S(n6768), .Z(n6358)
         );
  MUX2_X1 U6416 ( .A(n6358), .B(n6357), .S(n6731), .Z(n6359) );
  MUX2_X1 U6417 ( .A(n6359), .B(n6356), .S(n6714), .Z(n6360) );
  MUX2_X1 U6418 ( .A(n6360), .B(n6353), .S(n6705), .Z(n6361) );
  MUX2_X1 U6419 ( .A(reg_mem[1422]), .B(reg_mem[1414]), .S(n6769), .Z(n6362)
         );
  MUX2_X1 U6420 ( .A(reg_mem[1438]), .B(reg_mem[1430]), .S(n6769), .Z(n6363)
         );
  MUX2_X1 U6421 ( .A(n6363), .B(n6362), .S(n6732), .Z(n6364) );
  MUX2_X1 U6422 ( .A(reg_mem[1454]), .B(reg_mem[1446]), .S(n6769), .Z(n6365)
         );
  MUX2_X1 U6423 ( .A(reg_mem[1470]), .B(reg_mem[1462]), .S(n6769), .Z(n6366)
         );
  MUX2_X1 U6424 ( .A(n6366), .B(n6365), .S(n6732), .Z(n6367) );
  MUX2_X1 U6425 ( .A(n6367), .B(n6364), .S(n6714), .Z(n6368) );
  MUX2_X1 U6426 ( .A(reg_mem[1486]), .B(reg_mem[1478]), .S(n6769), .Z(n6369)
         );
  MUX2_X1 U6427 ( .A(reg_mem[1502]), .B(reg_mem[1494]), .S(n6769), .Z(n6370)
         );
  MUX2_X1 U6428 ( .A(n6370), .B(n6369), .S(n6732), .Z(n6371) );
  MUX2_X1 U6429 ( .A(reg_mem[1518]), .B(reg_mem[1510]), .S(n6769), .Z(n6372)
         );
  MUX2_X1 U6430 ( .A(reg_mem[1534]), .B(reg_mem[1526]), .S(n6769), .Z(n6373)
         );
  MUX2_X1 U6431 ( .A(n6373), .B(n6372), .S(n6732), .Z(n6374) );
  MUX2_X1 U6432 ( .A(n6374), .B(n6371), .S(n6714), .Z(n6375) );
  MUX2_X1 U6433 ( .A(n6375), .B(n6368), .S(n6705), .Z(n6376) );
  MUX2_X1 U6434 ( .A(n6376), .B(n6361), .S(n6699), .Z(n6377) );
  MUX2_X1 U6435 ( .A(n6377), .B(n6346), .S(n6697), .Z(n6378) );
  MUX2_X1 U6436 ( .A(reg_mem[1550]), .B(reg_mem[1542]), .S(n6769), .Z(n6379)
         );
  MUX2_X1 U6437 ( .A(reg_mem[1566]), .B(reg_mem[1558]), .S(n6769), .Z(n6380)
         );
  MUX2_X1 U6438 ( .A(n6380), .B(n6379), .S(n6732), .Z(n6381) );
  MUX2_X1 U6439 ( .A(reg_mem[1582]), .B(reg_mem[1574]), .S(n6769), .Z(n6382)
         );
  MUX2_X1 U6440 ( .A(reg_mem[1598]), .B(reg_mem[1590]), .S(n6769), .Z(n6383)
         );
  MUX2_X1 U6441 ( .A(n6383), .B(n6382), .S(n6732), .Z(n6384) );
  MUX2_X1 U6442 ( .A(n6384), .B(n6381), .S(n6714), .Z(n6385) );
  MUX2_X1 U6443 ( .A(reg_mem[1614]), .B(reg_mem[1606]), .S(n6770), .Z(n6386)
         );
  MUX2_X1 U6444 ( .A(reg_mem[1630]), .B(reg_mem[1622]), .S(n6770), .Z(n6387)
         );
  MUX2_X1 U6445 ( .A(n6387), .B(n6386), .S(n6732), .Z(n6388) );
  MUX2_X1 U6446 ( .A(reg_mem[1646]), .B(reg_mem[1638]), .S(n6770), .Z(n6389)
         );
  MUX2_X1 U6447 ( .A(reg_mem[1662]), .B(reg_mem[1654]), .S(n6770), .Z(n6390)
         );
  MUX2_X1 U6448 ( .A(n6390), .B(n6389), .S(n6732), .Z(n6391) );
  MUX2_X1 U6449 ( .A(n6391), .B(n6388), .S(n6714), .Z(n6392) );
  MUX2_X1 U6450 ( .A(n6392), .B(n6385), .S(n6705), .Z(n6393) );
  MUX2_X1 U6451 ( .A(reg_mem[1678]), .B(reg_mem[1670]), .S(n6770), .Z(n6394)
         );
  MUX2_X1 U6452 ( .A(reg_mem[1694]), .B(reg_mem[1686]), .S(n6770), .Z(n6395)
         );
  MUX2_X1 U6453 ( .A(n6395), .B(n6394), .S(n6732), .Z(n6396) );
  MUX2_X1 U6454 ( .A(reg_mem[1710]), .B(reg_mem[1702]), .S(n6770), .Z(n6397)
         );
  MUX2_X1 U6455 ( .A(reg_mem[1726]), .B(reg_mem[1718]), .S(n6770), .Z(n6398)
         );
  MUX2_X1 U6456 ( .A(n6398), .B(n6397), .S(n6732), .Z(n6399) );
  MUX2_X1 U6457 ( .A(n6399), .B(n6396), .S(n6714), .Z(n6400) );
  MUX2_X1 U6458 ( .A(reg_mem[1742]), .B(reg_mem[1734]), .S(n6770), .Z(n6401)
         );
  MUX2_X1 U6459 ( .A(reg_mem[1758]), .B(reg_mem[1750]), .S(n6770), .Z(n6402)
         );
  MUX2_X1 U6460 ( .A(n6402), .B(n6401), .S(n6732), .Z(n6403) );
  MUX2_X1 U6461 ( .A(reg_mem[1774]), .B(reg_mem[1766]), .S(n6770), .Z(n6404)
         );
  MUX2_X1 U6462 ( .A(reg_mem[1790]), .B(reg_mem[1782]), .S(n6770), .Z(n6405)
         );
  MUX2_X1 U6463 ( .A(n6405), .B(n6404), .S(n6732), .Z(n6406) );
  MUX2_X1 U6464 ( .A(n6406), .B(n6403), .S(n6714), .Z(n6407) );
  MUX2_X1 U6465 ( .A(n6407), .B(n6400), .S(n6705), .Z(n6408) );
  MUX2_X1 U6466 ( .A(n6408), .B(n6393), .S(n6699), .Z(n6409) );
  MUX2_X1 U6467 ( .A(reg_mem[1806]), .B(reg_mem[1798]), .S(n6771), .Z(n6410)
         );
  MUX2_X1 U6468 ( .A(reg_mem[1822]), .B(reg_mem[1814]), .S(n6771), .Z(n6411)
         );
  MUX2_X1 U6469 ( .A(n6411), .B(n6410), .S(n6733), .Z(n6412) );
  MUX2_X1 U6470 ( .A(reg_mem[1838]), .B(reg_mem[1830]), .S(n6771), .Z(n6413)
         );
  MUX2_X1 U6471 ( .A(reg_mem[1854]), .B(reg_mem[1846]), .S(n6771), .Z(n6414)
         );
  MUX2_X1 U6472 ( .A(n6414), .B(n6413), .S(n6733), .Z(n6415) );
  MUX2_X1 U6473 ( .A(n6415), .B(n6412), .S(n6715), .Z(n6416) );
  MUX2_X1 U6474 ( .A(reg_mem[1870]), .B(reg_mem[1862]), .S(n6771), .Z(n6417)
         );
  MUX2_X1 U6475 ( .A(reg_mem[1886]), .B(reg_mem[1878]), .S(n6771), .Z(n6418)
         );
  MUX2_X1 U6476 ( .A(n6418), .B(n6417), .S(n6733), .Z(n6419) );
  MUX2_X1 U6477 ( .A(reg_mem[1902]), .B(reg_mem[1894]), .S(n6771), .Z(n6420)
         );
  MUX2_X1 U6478 ( .A(reg_mem[1918]), .B(reg_mem[1910]), .S(n6771), .Z(n6421)
         );
  MUX2_X1 U6479 ( .A(n6421), .B(n6420), .S(n6733), .Z(n6422) );
  MUX2_X1 U6480 ( .A(n6422), .B(n6419), .S(n6715), .Z(n6423) );
  MUX2_X1 U6481 ( .A(n6423), .B(n6416), .S(n6705), .Z(n6424) );
  MUX2_X1 U6482 ( .A(reg_mem[1934]), .B(reg_mem[1926]), .S(n6771), .Z(n6425)
         );
  MUX2_X1 U6483 ( .A(reg_mem[1950]), .B(reg_mem[1942]), .S(n6771), .Z(n6426)
         );
  MUX2_X1 U6484 ( .A(n6426), .B(n6425), .S(n6733), .Z(n6427) );
  MUX2_X1 U6485 ( .A(reg_mem[1966]), .B(reg_mem[1958]), .S(n6771), .Z(n6428)
         );
  MUX2_X1 U6486 ( .A(reg_mem[1982]), .B(reg_mem[1974]), .S(n6771), .Z(n6429)
         );
  MUX2_X1 U6487 ( .A(n6429), .B(n6428), .S(n6733), .Z(n6430) );
  MUX2_X1 U6488 ( .A(n6430), .B(n6427), .S(n6715), .Z(n6431) );
  MUX2_X1 U6489 ( .A(reg_mem[1998]), .B(reg_mem[1990]), .S(n6772), .Z(n6432)
         );
  MUX2_X1 U6490 ( .A(reg_mem[2014]), .B(reg_mem[2006]), .S(n6772), .Z(n6433)
         );
  MUX2_X1 U6491 ( .A(n6433), .B(n6432), .S(n6733), .Z(n6434) );
  MUX2_X1 U6492 ( .A(reg_mem[2030]), .B(reg_mem[2022]), .S(n6772), .Z(n6435)
         );
  MUX2_X1 U6493 ( .A(reg_mem[2046]), .B(reg_mem[2038]), .S(n6772), .Z(n6436)
         );
  MUX2_X1 U6494 ( .A(n6436), .B(n6435), .S(n6733), .Z(n6437) );
  MUX2_X1 U6495 ( .A(n6437), .B(n6434), .S(n6715), .Z(n6438) );
  MUX2_X1 U6496 ( .A(n6438), .B(n6431), .S(n6705), .Z(n6439) );
  MUX2_X1 U6497 ( .A(n6439), .B(n6424), .S(n6699), .Z(n6440) );
  MUX2_X1 U6498 ( .A(n6440), .B(n6409), .S(n6697), .Z(n6441) );
  MUX2_X1 U6499 ( .A(n6441), .B(n6378), .S(addr_r[6]), .Z(n6442) );
  MUX2_X1 U6500 ( .A(n6442), .B(n6315), .S(addr_r[7]), .Z(data_r[6]) );
  MUX2_X1 U6501 ( .A(reg_mem[15]), .B(reg_mem[7]), .S(n6772), .Z(n6443) );
  MUX2_X1 U6502 ( .A(reg_mem[31]), .B(reg_mem[23]), .S(n6772), .Z(n6444) );
  MUX2_X1 U6503 ( .A(n6444), .B(n6443), .S(n6733), .Z(n6445) );
  MUX2_X1 U6504 ( .A(reg_mem[47]), .B(reg_mem[39]), .S(n6772), .Z(n6446) );
  MUX2_X1 U6505 ( .A(reg_mem[63]), .B(reg_mem[55]), .S(n6772), .Z(n6447) );
  MUX2_X1 U6506 ( .A(n6447), .B(n6446), .S(n6733), .Z(n6448) );
  MUX2_X1 U6507 ( .A(n6448), .B(n6445), .S(n6715), .Z(n6449) );
  MUX2_X1 U6508 ( .A(reg_mem[79]), .B(reg_mem[71]), .S(n6772), .Z(n6450) );
  MUX2_X1 U6509 ( .A(reg_mem[95]), .B(reg_mem[87]), .S(n6772), .Z(n6451) );
  MUX2_X1 U6510 ( .A(n6451), .B(n6450), .S(n6733), .Z(n6452) );
  MUX2_X1 U6511 ( .A(reg_mem[111]), .B(reg_mem[103]), .S(n6772), .Z(n6453) );
  MUX2_X1 U6512 ( .A(reg_mem[127]), .B(reg_mem[119]), .S(n6772), .Z(n6454) );
  MUX2_X1 U6513 ( .A(n6454), .B(n6453), .S(n6733), .Z(n6455) );
  MUX2_X1 U6514 ( .A(n6455), .B(n6452), .S(n6715), .Z(n6456) );
  MUX2_X1 U6515 ( .A(n6456), .B(n6449), .S(n6705), .Z(n6457) );
  MUX2_X1 U6516 ( .A(reg_mem[143]), .B(reg_mem[135]), .S(n6773), .Z(n6458) );
  MUX2_X1 U6517 ( .A(reg_mem[159]), .B(reg_mem[151]), .S(n6773), .Z(n6459) );
  MUX2_X1 U6518 ( .A(n6459), .B(n6458), .S(n6734), .Z(n6460) );
  MUX2_X1 U6519 ( .A(reg_mem[175]), .B(reg_mem[167]), .S(n6773), .Z(n6461) );
  MUX2_X1 U6520 ( .A(reg_mem[191]), .B(reg_mem[183]), .S(n6773), .Z(n6462) );
  MUX2_X1 U6521 ( .A(n6462), .B(n6461), .S(n6734), .Z(n6463) );
  MUX2_X1 U6522 ( .A(n6463), .B(n6460), .S(n6715), .Z(n6464) );
  MUX2_X1 U6523 ( .A(reg_mem[207]), .B(reg_mem[199]), .S(n6773), .Z(n6465) );
  MUX2_X1 U6524 ( .A(reg_mem[223]), .B(reg_mem[215]), .S(n6773), .Z(n6466) );
  MUX2_X1 U6525 ( .A(n6466), .B(n6465), .S(n6734), .Z(n6467) );
  MUX2_X1 U6526 ( .A(reg_mem[239]), .B(reg_mem[231]), .S(n6773), .Z(n6468) );
  MUX2_X1 U6527 ( .A(reg_mem[255]), .B(reg_mem[247]), .S(n6773), .Z(n6469) );
  MUX2_X1 U6528 ( .A(n6469), .B(n6468), .S(n6734), .Z(n6470) );
  MUX2_X1 U6529 ( .A(n6470), .B(n6467), .S(n6715), .Z(n6471) );
  MUX2_X1 U6530 ( .A(n6471), .B(n6464), .S(n6705), .Z(n6472) );
  MUX2_X1 U6531 ( .A(n6472), .B(n6457), .S(n6699), .Z(n6473) );
  MUX2_X1 U6532 ( .A(reg_mem[271]), .B(reg_mem[263]), .S(n6773), .Z(n6474) );
  MUX2_X1 U6533 ( .A(reg_mem[287]), .B(reg_mem[279]), .S(n6773), .Z(n6475) );
  MUX2_X1 U6534 ( .A(n6475), .B(n6474), .S(n6734), .Z(n6476) );
  MUX2_X1 U6535 ( .A(reg_mem[303]), .B(reg_mem[295]), .S(n6773), .Z(n6477) );
  MUX2_X1 U6536 ( .A(reg_mem[319]), .B(reg_mem[311]), .S(n6773), .Z(n6478) );
  MUX2_X1 U6537 ( .A(n6478), .B(n6477), .S(n6734), .Z(n6479) );
  MUX2_X1 U6538 ( .A(n6479), .B(n6476), .S(n6715), .Z(n6480) );
  MUX2_X1 U6539 ( .A(reg_mem[335]), .B(reg_mem[327]), .S(n6774), .Z(n6481) );
  MUX2_X1 U6540 ( .A(reg_mem[351]), .B(reg_mem[343]), .S(n6774), .Z(n6482) );
  MUX2_X1 U6541 ( .A(n6482), .B(n6481), .S(n6734), .Z(n6483) );
  MUX2_X1 U6542 ( .A(reg_mem[367]), .B(reg_mem[359]), .S(n6774), .Z(n6484) );
  MUX2_X1 U6543 ( .A(reg_mem[383]), .B(reg_mem[375]), .S(n6774), .Z(n6485) );
  MUX2_X1 U6544 ( .A(n6485), .B(n6484), .S(n6734), .Z(n6486) );
  MUX2_X1 U6545 ( .A(n6486), .B(n6483), .S(n6715), .Z(n6487) );
  MUX2_X1 U6546 ( .A(n6487), .B(n6480), .S(n6705), .Z(n6488) );
  MUX2_X1 U6547 ( .A(reg_mem[399]), .B(reg_mem[391]), .S(n6774), .Z(n6489) );
  MUX2_X1 U6548 ( .A(reg_mem[415]), .B(reg_mem[407]), .S(n6774), .Z(n6490) );
  MUX2_X1 U6549 ( .A(n6490), .B(n6489), .S(n6734), .Z(n6491) );
  MUX2_X1 U6550 ( .A(reg_mem[431]), .B(reg_mem[423]), .S(n6774), .Z(n6492) );
  MUX2_X1 U6551 ( .A(reg_mem[447]), .B(reg_mem[439]), .S(n6774), .Z(n6493) );
  MUX2_X1 U6552 ( .A(n6493), .B(n6492), .S(n6734), .Z(n6494) );
  MUX2_X1 U6553 ( .A(n6494), .B(n6491), .S(n6715), .Z(n6495) );
  MUX2_X1 U6554 ( .A(reg_mem[463]), .B(reg_mem[455]), .S(n6774), .Z(n6496) );
  MUX2_X1 U6555 ( .A(reg_mem[479]), .B(reg_mem[471]), .S(n6774), .Z(n6497) );
  MUX2_X1 U6556 ( .A(n6497), .B(n6496), .S(n6734), .Z(n6498) );
  MUX2_X1 U6557 ( .A(reg_mem[495]), .B(reg_mem[487]), .S(n6774), .Z(n6499) );
  MUX2_X1 U6558 ( .A(reg_mem[511]), .B(reg_mem[503]), .S(n6774), .Z(n6500) );
  MUX2_X1 U6559 ( .A(n6500), .B(n6499), .S(n6734), .Z(n6501) );
  MUX2_X1 U6560 ( .A(n6501), .B(n6498), .S(n6715), .Z(n6502) );
  MUX2_X1 U6561 ( .A(n6502), .B(n6495), .S(n6705), .Z(n6503) );
  MUX2_X1 U6562 ( .A(n6503), .B(n6488), .S(n6699), .Z(n6504) );
  MUX2_X1 U6563 ( .A(n6504), .B(n6473), .S(n6697), .Z(n6505) );
  MUX2_X1 U6564 ( .A(reg_mem[527]), .B(reg_mem[519]), .S(n6775), .Z(n6506) );
  MUX2_X1 U6565 ( .A(reg_mem[543]), .B(reg_mem[535]), .S(n6775), .Z(n6507) );
  MUX2_X1 U6566 ( .A(n6507), .B(n6506), .S(n6735), .Z(n6508) );
  MUX2_X1 U6567 ( .A(reg_mem[559]), .B(reg_mem[551]), .S(n6775), .Z(n6509) );
  MUX2_X1 U6568 ( .A(reg_mem[575]), .B(reg_mem[567]), .S(n6775), .Z(n6510) );
  MUX2_X1 U6569 ( .A(n6510), .B(n6509), .S(n6735), .Z(n6511) );
  MUX2_X1 U6570 ( .A(n6511), .B(n6508), .S(n6713), .Z(n6512) );
  MUX2_X1 U6571 ( .A(reg_mem[591]), .B(reg_mem[583]), .S(n6775), .Z(n6513) );
  MUX2_X1 U6572 ( .A(reg_mem[607]), .B(reg_mem[599]), .S(n6775), .Z(n6514) );
  MUX2_X1 U6573 ( .A(n6514), .B(n6513), .S(n6735), .Z(n6515) );
  MUX2_X1 U6574 ( .A(reg_mem[623]), .B(reg_mem[615]), .S(n6775), .Z(n6516) );
  MUX2_X1 U6575 ( .A(reg_mem[639]), .B(reg_mem[631]), .S(n6775), .Z(n6517) );
  MUX2_X1 U6576 ( .A(n6517), .B(n6516), .S(n6735), .Z(n6518) );
  MUX2_X1 U6577 ( .A(n6518), .B(n6515), .S(n6712), .Z(n6519) );
  MUX2_X1 U6578 ( .A(n6519), .B(n6512), .S(n6706), .Z(n6520) );
  MUX2_X1 U6579 ( .A(reg_mem[655]), .B(reg_mem[647]), .S(n6775), .Z(n6521) );
  MUX2_X1 U6580 ( .A(reg_mem[671]), .B(reg_mem[663]), .S(n6775), .Z(n6522) );
  MUX2_X1 U6581 ( .A(n6522), .B(n6521), .S(n6735), .Z(n6523) );
  MUX2_X1 U6582 ( .A(reg_mem[687]), .B(reg_mem[679]), .S(n6775), .Z(n6524) );
  MUX2_X1 U6583 ( .A(reg_mem[703]), .B(reg_mem[695]), .S(n6775), .Z(n6525) );
  MUX2_X1 U6584 ( .A(n6525), .B(n6524), .S(n6735), .Z(n6526) );
  MUX2_X1 U6585 ( .A(n6526), .B(n6523), .S(n6709), .Z(n6527) );
  MUX2_X1 U6586 ( .A(reg_mem[719]), .B(reg_mem[711]), .S(n6776), .Z(n6528) );
  MUX2_X1 U6587 ( .A(reg_mem[735]), .B(reg_mem[727]), .S(n6776), .Z(n6529) );
  MUX2_X1 U6588 ( .A(n6529), .B(n6528), .S(n6735), .Z(n6530) );
  MUX2_X1 U6589 ( .A(reg_mem[751]), .B(reg_mem[743]), .S(n6776), .Z(n6531) );
  MUX2_X1 U6590 ( .A(reg_mem[767]), .B(reg_mem[759]), .S(n6776), .Z(n6532) );
  MUX2_X1 U6591 ( .A(n6532), .B(n6531), .S(n6735), .Z(n6533) );
  MUX2_X1 U6592 ( .A(n6533), .B(n6530), .S(n6717), .Z(n6534) );
  MUX2_X1 U6593 ( .A(n6534), .B(n6527), .S(n6706), .Z(n6535) );
  MUX2_X1 U6594 ( .A(n6535), .B(n6520), .S(n6699), .Z(n6536) );
  MUX2_X1 U6595 ( .A(reg_mem[783]), .B(reg_mem[775]), .S(n6776), .Z(n6537) );
  MUX2_X1 U6596 ( .A(reg_mem[799]), .B(reg_mem[791]), .S(n6776), .Z(n6538) );
  MUX2_X1 U6597 ( .A(n6538), .B(n6537), .S(n6735), .Z(n6539) );
  MUX2_X1 U6598 ( .A(reg_mem[815]), .B(reg_mem[807]), .S(n6776), .Z(n6540) );
  MUX2_X1 U6599 ( .A(reg_mem[831]), .B(reg_mem[823]), .S(n6776), .Z(n6541) );
  MUX2_X1 U6600 ( .A(n6541), .B(n6540), .S(n6735), .Z(n6542) );
  MUX2_X1 U6601 ( .A(n6542), .B(n6539), .S(n6715), .Z(n6543) );
  MUX2_X1 U6602 ( .A(reg_mem[847]), .B(reg_mem[839]), .S(n6776), .Z(n6544) );
  MUX2_X1 U6603 ( .A(reg_mem[863]), .B(reg_mem[855]), .S(n6776), .Z(n6545) );
  MUX2_X1 U6604 ( .A(n6545), .B(n6544), .S(n6735), .Z(n6546) );
  MUX2_X1 U6605 ( .A(reg_mem[879]), .B(reg_mem[871]), .S(n6776), .Z(n6547) );
  MUX2_X1 U6606 ( .A(reg_mem[895]), .B(reg_mem[887]), .S(n6776), .Z(n6548) );
  MUX2_X1 U6607 ( .A(n6548), .B(n6547), .S(n6735), .Z(n6549) );
  MUX2_X1 U6608 ( .A(n6549), .B(n6546), .S(n6711), .Z(n6550) );
  MUX2_X1 U6609 ( .A(n6550), .B(n6543), .S(n6706), .Z(n6551) );
  MUX2_X1 U6610 ( .A(reg_mem[911]), .B(reg_mem[903]), .S(n6777), .Z(n6552) );
  MUX2_X1 U6611 ( .A(reg_mem[927]), .B(reg_mem[919]), .S(n6777), .Z(n6553) );
  MUX2_X1 U6612 ( .A(n6553), .B(n6552), .S(n6736), .Z(n6554) );
  MUX2_X1 U6613 ( .A(reg_mem[943]), .B(reg_mem[935]), .S(n6777), .Z(n6555) );
  MUX2_X1 U6614 ( .A(reg_mem[959]), .B(reg_mem[951]), .S(n6777), .Z(n6556) );
  MUX2_X1 U6615 ( .A(n6556), .B(n6555), .S(n6736), .Z(n6557) );
  MUX2_X1 U6616 ( .A(n6557), .B(n6554), .S(n6707), .Z(n6558) );
  MUX2_X1 U6617 ( .A(reg_mem[975]), .B(reg_mem[967]), .S(n6777), .Z(n6559) );
  MUX2_X1 U6618 ( .A(reg_mem[991]), .B(reg_mem[983]), .S(n6777), .Z(n6560) );
  MUX2_X1 U6619 ( .A(n6560), .B(n6559), .S(n6736), .Z(n6561) );
  MUX2_X1 U6620 ( .A(reg_mem[1007]), .B(reg_mem[999]), .S(n6777), .Z(n6562) );
  MUX2_X1 U6621 ( .A(reg_mem[1023]), .B(reg_mem[1015]), .S(n6777), .Z(n6563)
         );
  MUX2_X1 U6622 ( .A(n6563), .B(n6562), .S(n6736), .Z(n6564) );
  MUX2_X1 U6623 ( .A(n6564), .B(n6561), .S(n6713), .Z(n6565) );
  MUX2_X1 U6624 ( .A(n6565), .B(n6558), .S(n6706), .Z(n6566) );
  MUX2_X1 U6625 ( .A(n6566), .B(n6551), .S(n6699), .Z(n6567) );
  MUX2_X1 U6626 ( .A(n6567), .B(n6536), .S(n6697), .Z(n6568) );
  MUX2_X1 U6627 ( .A(n6568), .B(n6505), .S(addr_r[6]), .Z(n6569) );
  MUX2_X1 U6628 ( .A(reg_mem[1039]), .B(reg_mem[1031]), .S(n6777), .Z(n6570)
         );
  MUX2_X1 U6629 ( .A(reg_mem[1055]), .B(reg_mem[1047]), .S(n6777), .Z(n6571)
         );
  MUX2_X1 U6630 ( .A(n6571), .B(n6570), .S(n6736), .Z(n6572) );
  MUX2_X1 U6631 ( .A(reg_mem[1071]), .B(reg_mem[1063]), .S(n6777), .Z(n6573)
         );
  MUX2_X1 U6632 ( .A(reg_mem[1087]), .B(reg_mem[1079]), .S(n6777), .Z(n6574)
         );
  MUX2_X1 U6633 ( .A(n6574), .B(n6573), .S(n6736), .Z(n6575) );
  MUX2_X1 U6634 ( .A(n6575), .B(n6572), .S(n6710), .Z(n6576) );
  MUX2_X1 U6635 ( .A(reg_mem[1103]), .B(reg_mem[1095]), .S(n6778), .Z(n6577)
         );
  MUX2_X1 U6636 ( .A(reg_mem[1119]), .B(reg_mem[1111]), .S(n6778), .Z(n6578)
         );
  MUX2_X1 U6637 ( .A(n6578), .B(n6577), .S(n6736), .Z(n6579) );
  MUX2_X1 U6638 ( .A(reg_mem[1135]), .B(reg_mem[1127]), .S(n6778), .Z(n6580)
         );
  MUX2_X1 U6639 ( .A(reg_mem[1151]), .B(reg_mem[1143]), .S(n6778), .Z(n6581)
         );
  MUX2_X1 U6640 ( .A(n6581), .B(n6580), .S(n6736), .Z(n6582) );
  MUX2_X1 U6641 ( .A(n6582), .B(n6579), .S(n6716), .Z(n6583) );
  MUX2_X1 U6642 ( .A(n6583), .B(n6576), .S(n6706), .Z(n6584) );
  MUX2_X1 U6643 ( .A(reg_mem[1167]), .B(reg_mem[1159]), .S(n6778), .Z(n6585)
         );
  MUX2_X1 U6644 ( .A(reg_mem[1183]), .B(reg_mem[1175]), .S(n6778), .Z(n6586)
         );
  MUX2_X1 U6645 ( .A(n6586), .B(n6585), .S(n6736), .Z(n6587) );
  MUX2_X1 U6646 ( .A(reg_mem[1199]), .B(reg_mem[1191]), .S(n6778), .Z(n6588)
         );
  MUX2_X1 U6647 ( .A(reg_mem[1215]), .B(reg_mem[1207]), .S(n6778), .Z(n6589)
         );
  MUX2_X1 U6648 ( .A(n6589), .B(n6588), .S(n6736), .Z(n6590) );
  MUX2_X1 U6649 ( .A(n6590), .B(n6587), .S(n6708), .Z(n6591) );
  MUX2_X1 U6650 ( .A(reg_mem[1231]), .B(reg_mem[1223]), .S(n6778), .Z(n6592)
         );
  MUX2_X1 U6651 ( .A(reg_mem[1247]), .B(reg_mem[1239]), .S(n6778), .Z(n6593)
         );
  MUX2_X1 U6652 ( .A(n6593), .B(n6592), .S(n6736), .Z(n6594) );
  MUX2_X1 U6653 ( .A(reg_mem[1263]), .B(reg_mem[1255]), .S(n6778), .Z(n6595)
         );
  MUX2_X1 U6654 ( .A(reg_mem[1279]), .B(reg_mem[1271]), .S(n6778), .Z(n6596)
         );
  MUX2_X1 U6655 ( .A(n6596), .B(n6595), .S(n6736), .Z(n6597) );
  MUX2_X1 U6656 ( .A(n6597), .B(n6594), .S(n6714), .Z(n6598) );
  MUX2_X1 U6657 ( .A(n6598), .B(n6591), .S(n6706), .Z(n6599) );
  MUX2_X1 U6658 ( .A(n6599), .B(n6584), .S(n6699), .Z(n6600) );
  MUX2_X1 U6659 ( .A(reg_mem[1295]), .B(reg_mem[1287]), .S(n6779), .Z(n6601)
         );
  MUX2_X1 U6660 ( .A(reg_mem[1311]), .B(reg_mem[1303]), .S(n6779), .Z(n6602)
         );
  MUX2_X1 U6661 ( .A(n6602), .B(n6601), .S(n6737), .Z(n6603) );
  MUX2_X1 U6662 ( .A(reg_mem[1327]), .B(reg_mem[1319]), .S(n6779), .Z(n6604)
         );
  MUX2_X1 U6663 ( .A(reg_mem[1343]), .B(reg_mem[1335]), .S(n6779), .Z(n6605)
         );
  MUX2_X1 U6664 ( .A(n6605), .B(n6604), .S(n6737), .Z(n6606) );
  MUX2_X1 U6665 ( .A(n6606), .B(n6603), .S(n6716), .Z(n6607) );
  MUX2_X1 U6666 ( .A(reg_mem[1359]), .B(reg_mem[1351]), .S(n6779), .Z(n6608)
         );
  MUX2_X1 U6667 ( .A(reg_mem[1375]), .B(reg_mem[1367]), .S(n6779), .Z(n6609)
         );
  MUX2_X1 U6668 ( .A(n6609), .B(n6608), .S(n6737), .Z(n6610) );
  MUX2_X1 U6669 ( .A(reg_mem[1391]), .B(reg_mem[1383]), .S(n6779), .Z(n6611)
         );
  MUX2_X1 U6670 ( .A(reg_mem[1407]), .B(reg_mem[1399]), .S(n6779), .Z(n6612)
         );
  MUX2_X1 U6671 ( .A(n6612), .B(n6611), .S(n6737), .Z(n6613) );
  MUX2_X1 U6672 ( .A(n6613), .B(n6610), .S(n6716), .Z(n6614) );
  MUX2_X1 U6673 ( .A(n6614), .B(n6607), .S(n6706), .Z(n6615) );
  MUX2_X1 U6674 ( .A(reg_mem[1423]), .B(reg_mem[1415]), .S(n6779), .Z(n6616)
         );
  MUX2_X1 U6675 ( .A(reg_mem[1439]), .B(reg_mem[1431]), .S(n6779), .Z(n6617)
         );
  MUX2_X1 U6676 ( .A(n6617), .B(n6616), .S(n6737), .Z(n6618) );
  MUX2_X1 U6677 ( .A(reg_mem[1455]), .B(reg_mem[1447]), .S(n6779), .Z(n6619)
         );
  MUX2_X1 U6678 ( .A(reg_mem[1471]), .B(reg_mem[1463]), .S(n6779), .Z(n6620)
         );
  MUX2_X1 U6679 ( .A(n6620), .B(n6619), .S(n6737), .Z(n6621) );
  MUX2_X1 U6680 ( .A(n6621), .B(n6618), .S(n6716), .Z(n6622) );
  MUX2_X1 U6681 ( .A(reg_mem[1487]), .B(reg_mem[1479]), .S(n6780), .Z(n6623)
         );
  MUX2_X1 U6682 ( .A(reg_mem[1503]), .B(reg_mem[1495]), .S(n6780), .Z(n6624)
         );
  MUX2_X1 U6683 ( .A(n6624), .B(n6623), .S(n6737), .Z(n6625) );
  MUX2_X1 U6684 ( .A(reg_mem[1519]), .B(reg_mem[1511]), .S(n6780), .Z(n6626)
         );
  MUX2_X1 U6685 ( .A(reg_mem[1535]), .B(reg_mem[1527]), .S(n6780), .Z(n6627)
         );
  MUX2_X1 U6686 ( .A(n6627), .B(n6626), .S(n6737), .Z(n6628) );
  MUX2_X1 U6687 ( .A(n6628), .B(n6625), .S(n6716), .Z(n6629) );
  MUX2_X1 U6688 ( .A(n6629), .B(n6622), .S(n6706), .Z(n6630) );
  MUX2_X1 U6689 ( .A(n6630), .B(n6615), .S(n6699), .Z(n6631) );
  MUX2_X1 U6690 ( .A(n6631), .B(n6600), .S(n6697), .Z(n6632) );
  MUX2_X1 U6691 ( .A(reg_mem[1551]), .B(reg_mem[1543]), .S(n6780), .Z(n6633)
         );
  MUX2_X1 U6692 ( .A(reg_mem[1567]), .B(reg_mem[1559]), .S(n6780), .Z(n6634)
         );
  MUX2_X1 U6693 ( .A(n6634), .B(n6633), .S(n6737), .Z(n6635) );
  MUX2_X1 U6694 ( .A(reg_mem[1583]), .B(reg_mem[1575]), .S(n6780), .Z(n6636)
         );
  MUX2_X1 U6695 ( .A(reg_mem[1599]), .B(reg_mem[1591]), .S(n6780), .Z(n6637)
         );
  MUX2_X1 U6696 ( .A(n6637), .B(n6636), .S(n6737), .Z(n6638) );
  MUX2_X1 U6697 ( .A(n6638), .B(n6635), .S(n6716), .Z(n6639) );
  MUX2_X1 U6698 ( .A(reg_mem[1615]), .B(reg_mem[1607]), .S(n6780), .Z(n6640)
         );
  MUX2_X1 U6699 ( .A(reg_mem[1631]), .B(reg_mem[1623]), .S(n6780), .Z(n6641)
         );
  MUX2_X1 U6700 ( .A(n6641), .B(n6640), .S(n6737), .Z(n6642) );
  MUX2_X1 U6701 ( .A(reg_mem[1647]), .B(reg_mem[1639]), .S(n6780), .Z(n6643)
         );
  MUX2_X1 U6702 ( .A(reg_mem[1663]), .B(reg_mem[1655]), .S(n6780), .Z(n6644)
         );
  MUX2_X1 U6703 ( .A(n6644), .B(n6643), .S(n6737), .Z(n6645) );
  MUX2_X1 U6704 ( .A(n6645), .B(n6642), .S(n6716), .Z(n6646) );
  MUX2_X1 U6705 ( .A(n6646), .B(n6639), .S(n6706), .Z(n6647) );
  MUX2_X1 U6706 ( .A(reg_mem[1679]), .B(reg_mem[1671]), .S(n6781), .Z(n6648)
         );
  MUX2_X1 U6707 ( .A(reg_mem[1695]), .B(reg_mem[1687]), .S(n6781), .Z(n6649)
         );
  MUX2_X1 U6708 ( .A(n6649), .B(n6648), .S(n6738), .Z(n6650) );
  MUX2_X1 U6709 ( .A(reg_mem[1711]), .B(reg_mem[1703]), .S(n6781), .Z(n6651)
         );
  MUX2_X1 U6710 ( .A(reg_mem[1727]), .B(reg_mem[1719]), .S(n6781), .Z(n6652)
         );
  MUX2_X1 U6711 ( .A(n6652), .B(n6651), .S(n6738), .Z(n6653) );
  MUX2_X1 U6712 ( .A(n6653), .B(n6650), .S(n6716), .Z(n6654) );
  MUX2_X1 U6713 ( .A(reg_mem[1743]), .B(reg_mem[1735]), .S(n6781), .Z(n6655)
         );
  MUX2_X1 U6714 ( .A(reg_mem[1759]), .B(reg_mem[1751]), .S(n6781), .Z(n6656)
         );
  MUX2_X1 U6715 ( .A(n6656), .B(n6655), .S(n6738), .Z(n6657) );
  MUX2_X1 U6716 ( .A(reg_mem[1775]), .B(reg_mem[1767]), .S(n6781), .Z(n6658)
         );
  MUX2_X1 U6717 ( .A(reg_mem[1791]), .B(reg_mem[1783]), .S(n6781), .Z(n6659)
         );
  MUX2_X1 U6718 ( .A(n6659), .B(n6658), .S(n6738), .Z(n6660) );
  MUX2_X1 U6719 ( .A(n6660), .B(n6657), .S(n6716), .Z(n6661) );
  MUX2_X1 U6720 ( .A(n6661), .B(n6654), .S(n6706), .Z(n6662) );
  MUX2_X1 U6721 ( .A(n6662), .B(n6647), .S(n6699), .Z(n6663) );
  MUX2_X1 U6722 ( .A(reg_mem[1807]), .B(reg_mem[1799]), .S(n6781), .Z(n6664)
         );
  MUX2_X1 U6723 ( .A(reg_mem[1823]), .B(reg_mem[1815]), .S(n6781), .Z(n6665)
         );
  MUX2_X1 U6724 ( .A(n6665), .B(n6664), .S(n6738), .Z(n6666) );
  MUX2_X1 U6725 ( .A(reg_mem[1839]), .B(reg_mem[1831]), .S(n6781), .Z(n6667)
         );
  MUX2_X1 U6726 ( .A(reg_mem[1855]), .B(reg_mem[1847]), .S(n6781), .Z(n6668)
         );
  MUX2_X1 U6727 ( .A(n6668), .B(n6667), .S(n6738), .Z(n6669) );
  MUX2_X1 U6728 ( .A(n6669), .B(n6666), .S(n6716), .Z(n6670) );
  MUX2_X1 U6729 ( .A(reg_mem[1871]), .B(reg_mem[1863]), .S(n6782), .Z(n6671)
         );
  MUX2_X1 U6730 ( .A(reg_mem[1887]), .B(reg_mem[1879]), .S(n6782), .Z(n6672)
         );
  MUX2_X1 U6731 ( .A(n6672), .B(n6671), .S(n6738), .Z(n6673) );
  MUX2_X1 U6732 ( .A(reg_mem[1903]), .B(reg_mem[1895]), .S(n6782), .Z(n6674)
         );
  MUX2_X1 U6733 ( .A(reg_mem[1919]), .B(reg_mem[1911]), .S(n6782), .Z(n6675)
         );
  MUX2_X1 U6734 ( .A(n6675), .B(n6674), .S(n6738), .Z(n6676) );
  MUX2_X1 U6735 ( .A(n6676), .B(n6673), .S(n6716), .Z(n6677) );
  MUX2_X1 U6736 ( .A(n6677), .B(n6670), .S(n6706), .Z(n6678) );
  MUX2_X1 U6737 ( .A(reg_mem[1935]), .B(reg_mem[1927]), .S(n6782), .Z(n6679)
         );
  MUX2_X1 U6738 ( .A(reg_mem[1951]), .B(reg_mem[1943]), .S(n6782), .Z(n6680)
         );
  MUX2_X1 U6739 ( .A(n6680), .B(n6679), .S(n6738), .Z(n6681) );
  MUX2_X1 U6740 ( .A(reg_mem[1967]), .B(reg_mem[1959]), .S(n6782), .Z(n6682)
         );
  MUX2_X1 U6741 ( .A(reg_mem[1983]), .B(reg_mem[1975]), .S(n6782), .Z(n6683)
         );
  MUX2_X1 U6742 ( .A(n6683), .B(n6682), .S(n6738), .Z(n6684) );
  MUX2_X1 U6743 ( .A(n6684), .B(n6681), .S(n6716), .Z(n6685) );
  MUX2_X1 U6744 ( .A(reg_mem[1999]), .B(reg_mem[1991]), .S(n6782), .Z(n6686)
         );
  MUX2_X1 U6745 ( .A(reg_mem[2015]), .B(reg_mem[2007]), .S(n6782), .Z(n6687)
         );
  MUX2_X1 U6746 ( .A(n6687), .B(n6686), .S(n6738), .Z(n6688) );
  MUX2_X1 U6747 ( .A(reg_mem[2031]), .B(reg_mem[2023]), .S(n6782), .Z(n6689)
         );
  MUX2_X1 U6748 ( .A(reg_mem[2047]), .B(reg_mem[2039]), .S(n6782), .Z(n6690)
         );
  MUX2_X1 U6749 ( .A(n6690), .B(n6689), .S(n6738), .Z(n6691) );
  MUX2_X1 U6750 ( .A(n6691), .B(n6688), .S(n6716), .Z(n6692) );
  MUX2_X1 U6751 ( .A(n6692), .B(n6685), .S(n6706), .Z(n6693) );
  MUX2_X1 U6752 ( .A(n6693), .B(n6678), .S(n6699), .Z(n6694) );
  MUX2_X1 U6753 ( .A(n6694), .B(n6663), .S(n6697), .Z(n6695) );
  MUX2_X1 U6754 ( .A(n6695), .B(n6632), .S(addr_r[6]), .Z(n6696) );
  MUX2_X1 U6755 ( .A(n6696), .B(n6569), .S(addr_r[7]), .Z(data_r[7]) );
  BUF_X1 U6756 ( .A(addr_r[4]), .Z(n6700) );
  BUF_X1 U6757 ( .A(addr_r[3]), .Z(n6702) );
  BUF_X1 U6758 ( .A(addr_r[3]), .Z(n6703) );
  BUF_X1 U6759 ( .A(addr_r[3]), .Z(n6704) );
  BUF_X1 U6760 ( .A(addr_r[3]), .Z(n6705) );
  BUF_X1 U6761 ( .A(addr_r[3]), .Z(n6706) );
  BUF_X1 U6762 ( .A(n6717), .Z(n6711) );
  BUF_X1 U6763 ( .A(n6717), .Z(n6712) );
  BUF_X1 U6764 ( .A(n6717), .Z(n6713) );
  BUF_X1 U6765 ( .A(n6717), .Z(n6714) );
  BUF_X1 U6766 ( .A(n6717), .Z(n6715) );
  BUF_X1 U6767 ( .A(n6717), .Z(n6716) );
  BUF_X1 U6768 ( .A(n6783), .Z(n6746) );
  BUF_X1 U6769 ( .A(n6781), .Z(n6747) );
  BUF_X1 U6770 ( .A(n6775), .Z(n6748) );
  BUF_X1 U6771 ( .A(n6782), .Z(n6749) );
  BUF_X1 U6772 ( .A(n6776), .Z(n6750) );
  BUF_X1 U6773 ( .A(n6742), .Z(n6751) );
  BUF_X1 U6774 ( .A(n6742), .Z(n6756) );
  BUF_X1 U6775 ( .A(n6742), .Z(n6757) );
  BUF_X1 U6776 ( .A(n6742), .Z(n6758) );
  BUF_X1 U6777 ( .A(n6742), .Z(n6759) );
  BUF_X1 U6778 ( .A(n6742), .Z(n6760) );
  BUF_X1 U6779 ( .A(n6742), .Z(n6761) );
  BUF_X1 U6780 ( .A(n6742), .Z(n6762) );
  BUF_X1 U6781 ( .A(n6741), .Z(n6767) );
  BUF_X1 U6782 ( .A(n6741), .Z(n6768) );
  BUF_X1 U6783 ( .A(n6741), .Z(n6769) );
  BUF_X1 U6784 ( .A(n6741), .Z(n6770) );
  BUF_X1 U6785 ( .A(n6741), .Z(n6771) );
  BUF_X1 U6786 ( .A(n6741), .Z(n6772) );
  BUF_X1 U6787 ( .A(n6741), .Z(n6773) );
  BUF_X1 U6788 ( .A(n6740), .Z(n6778) );
  BUF_X1 U6789 ( .A(n6740), .Z(n6779) );
  BUF_X1 U6790 ( .A(n6740), .Z(n6780) );
  BUF_X1 U6791 ( .A(n6740), .Z(n6781) );
  BUF_X1 U6792 ( .A(n6740), .Z(n6782) );
endmodule


module asyn_fifo_top_word_width8_1 ( r_clk, w_clk, rd, wr, reset_n, data_in, 
        data_out, full, empty );
  input [7:0] data_in;
  output [7:0] data_out;
  input r_clk, w_clk, rd, wr, reset_n;
  output full, empty;
  wire   we_enable;
  wire   [7:0] addr_r;
  wire   [7:0] addr_w;

  fifo_control_unit_addr_size8_1 fifo_ctrl ( .reset_n(reset_n), .w_clk(w_clk), 
        .r_clk(r_clk), .rd(rd), .wr(wr), .addr_r(addr_r), .addr_w(addr_w), 
        .full(full), .empty(empty), .we_enable(we_enable) );
  reg_memory_file_addr_size8_word_width8_1 fifo_memory ( .we_s(we_enable), 
        .clk(w_clk), .addr_r(addr_r), .addr_w(addr_w), .data_w(data_in), 
        .data_r(data_out) );
endmodule


module rx_D_bits9_sb_tick16 ( clk, reset_n, rx, s_tick, data_out, rx_done, 
        rx_err, fr_err );
  output [7:0] data_out;
  input clk, reset_n, rx, s_tick;
  output rx_done, rx_err, fr_err;
  wire   U3_U3_DATA4_2, U3_U3_DATA3_0, U3_U3_DATA3_1, U3_U3_DATA3_2,
         U3_U3_DATA3_3, U27_DATA2_0, U27_DATA2_1, U22_DATA1_0, n1, n2, n3, n4,
         n5, n6, n7, n13, n18, n19, n24, n25, n26, n27, n28, n29, n30, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180;

  XOR2_X1 U80 ( .A(U22_DATA1_0), .B(rx), .Z(n35) );
  DFFR_X1 n_reg_reg_1_ ( .D(n83), .CK(clk), .RN(reset_n), .QN(n29) );
  DFFR_X1 n_reg_reg_0_ ( .D(n92), .CK(clk), .RN(reset_n), .QN(n30) );
  DFFR_X1 b_reg_reg_0_ ( .D(n82), .CK(clk), .RN(reset_n), .Q(data_out[0]) );
  DFFR_X1 parity_reg_reg ( .D(n171), .CK(clk), .RN(reset_n), .Q(U22_DATA1_0)
         );
  DFFR_X1 b_reg_reg_6_ ( .D(n76), .CK(clk), .RN(reset_n), .Q(data_out[6]), 
        .QN(n2) );
  DFFR_X1 b_reg_reg_5_ ( .D(n77), .CK(clk), .RN(reset_n), .Q(data_out[5]), 
        .QN(n3) );
  DFFR_X1 b_reg_reg_4_ ( .D(n78), .CK(clk), .RN(reset_n), .Q(data_out[4]), 
        .QN(n4) );
  DFFR_X1 b_reg_reg_3_ ( .D(n79), .CK(clk), .RN(reset_n), .Q(data_out[3]), 
        .QN(n5) );
  DFFR_X1 b_reg_reg_2_ ( .D(n80), .CK(clk), .RN(reset_n), .Q(data_out[2]), 
        .QN(n6) );
  DFFR_X1 b_reg_reg_1_ ( .D(n81), .CK(clk), .RN(reset_n), .Q(data_out[1]), 
        .QN(n7) );
  DFFR_X1 b_reg_reg_7_ ( .D(n75), .CK(clk), .RN(reset_n), .Q(data_out[7]), 
        .QN(n1) );
  DFFR_X1 n_reg_reg_3_ ( .D(n91), .CK(clk), .RN(reset_n), .Q(n166), .QN(n27)
         );
  DFFR_X1 n_reg_reg_2_ ( .D(n84), .CK(clk), .RN(reset_n), .Q(U3_U3_DATA4_2), 
        .QN(n28) );
  DFFR_X1 s_reg_reg_3_ ( .D(n89), .CK(clk), .RN(reset_n), .Q(U3_U3_DATA3_3), 
        .QN(n19) );
  DFFR_X1 s_reg_reg_2_ ( .D(n87), .CK(clk), .RN(reset_n), .Q(U3_U3_DATA3_2), 
        .QN(n24) );
  DFFR_X1 s_reg_reg_1_ ( .D(n86), .CK(clk), .RN(reset_n), .Q(U3_U3_DATA3_1), 
        .QN(n25) );
  DFFR_X1 s_reg_reg_0_ ( .D(n85), .CK(clk), .RN(reset_n), .Q(U3_U3_DATA3_0), 
        .QN(n26) );
  DFFR_X1 state_reg_reg_1_ ( .D(n90), .CK(clk), .RN(reset_n), .Q(U27_DATA2_1), 
        .QN(n13) );
  DFFR_X1 state_reg_reg_0_ ( .D(n88), .CK(clk), .RN(reset_n), .Q(U27_DATA2_0), 
        .QN(n18) );
  NOR4_X1 U3 ( .A1(n24), .A2(n25), .A3(n26), .A4(U3_U3_DATA3_3), .ZN(n62) );
  INV_X1 U4 ( .A(n41), .ZN(n170) );
  OR2_X1 U5 ( .A1(n73), .A2(n68), .ZN(n45) );
  INV_X1 U6 ( .A(n73), .ZN(n173) );
  NAND2_X1 U7 ( .A1(s_tick), .A2(n175), .ZN(n66) );
  NOR2_X1 U8 ( .A1(n172), .A2(n40), .ZN(n41) );
  INV_X1 U9 ( .A(n38), .ZN(n172) );
  OAI21_X1 U10 ( .B1(n178), .B2(n177), .A(s_tick), .ZN(n68) );
  NAND2_X1 U11 ( .A1(s_tick), .A2(n178), .ZN(n40) );
  NOR2_X1 U12 ( .A1(n59), .A2(n179), .ZN(n74) );
  NAND2_X1 U13 ( .A1(n178), .A2(n38), .ZN(n73) );
  AND4_X1 U14 ( .A1(n35), .A2(n178), .A3(n167), .A4(n56), .ZN(rx_err) );
  INV_X1 U15 ( .A(n66), .ZN(n167) );
  AND2_X1 U16 ( .A1(n180), .A2(rx_done), .ZN(fr_err) );
  NOR2_X1 U17 ( .A1(n66), .A2(n69), .ZN(rx_done) );
  AOI211_X1 U18 ( .C1(n176), .C2(n177), .A(n168), .B(n178), .ZN(n54) );
  INV_X1 U19 ( .A(n62), .ZN(n176) );
  OAI21_X1 U20 ( .B1(n179), .B2(n59), .A(n60), .ZN(n49) );
  INV_X1 U21 ( .A(n57), .ZN(n168) );
  INV_X1 U22 ( .A(n37), .ZN(n178) );
  INV_X1 U23 ( .A(n64), .ZN(n175) );
  OAI22_X1 U24 ( .A1(n175), .A2(n37), .B1(n62), .B2(n70), .ZN(n59) );
  NOR2_X1 U25 ( .A1(n64), .A2(n56), .ZN(n38) );
  XNOR2_X1 U26 ( .A(n51), .B(n52), .ZN(n46) );
  XNOR2_X1 U27 ( .A(n48), .B(n50), .ZN(n44) );
  INV_X1 U28 ( .A(n70), .ZN(n177) );
  NAND3_X1 U29 ( .A1(n37), .A2(n69), .A3(n70), .ZN(n39) );
  NAND2_X1 U30 ( .A1(n50), .A2(n48), .ZN(n51) );
  INV_X1 U31 ( .A(n69), .ZN(n179) );
  INV_X1 U32 ( .A(rx), .ZN(n180) );
  AOI211_X1 U33 ( .C1(rx), .C2(n177), .A(n68), .B(n59), .ZN(n43) );
  OAI21_X1 U34 ( .B1(n18), .B2(n66), .A(n169), .ZN(n57) );
  OAI221_X1 U35 ( .B1(n168), .B2(n53), .C1(n54), .C2(n18), .A(n55), .ZN(n88)
         );
  NAND2_X1 U36 ( .A1(n18), .A2(n13), .ZN(n53) );
  NAND4_X1 U37 ( .A1(n56), .A2(n178), .A3(n175), .A4(n57), .ZN(n55) );
  OAI21_X1 U38 ( .B1(rx), .B2(n39), .A(n40), .ZN(n36) );
  AND2_X1 U39 ( .A1(n60), .A2(n61), .ZN(n47) );
  NAND3_X1 U40 ( .A1(n177), .A2(rx), .A3(n62), .ZN(n61) );
  OAI22_X1 U41 ( .A1(n47), .A2(n26), .B1(n48), .B2(n49), .ZN(n85) );
  OAI22_X1 U42 ( .A1(n43), .A2(n30), .B1(n48), .B2(n45), .ZN(n92) );
  OAI22_X1 U43 ( .A1(n47), .A2(n19), .B1(n49), .B2(n58), .ZN(n89) );
  OAI22_X1 U44 ( .A1(n41), .A2(n1), .B1(n180), .B2(n170), .ZN(n75) );
  OAI22_X1 U45 ( .A1(n47), .A2(n25), .B1(n44), .B2(n49), .ZN(n86) );
  OAI22_X1 U46 ( .A1(n47), .A2(n24), .B1(n46), .B2(n49), .ZN(n87) );
  OAI22_X1 U47 ( .A1(n43), .A2(n27), .B1(n45), .B2(n58), .ZN(n91) );
  OAI22_X1 U48 ( .A1(n43), .A2(n29), .B1(n44), .B2(n45), .ZN(n83) );
  OAI22_X1 U49 ( .A1(n43), .A2(n28), .B1(n45), .B2(n46), .ZN(n84) );
  OAI21_X1 U50 ( .B1(n54), .B2(n13), .A(n65), .ZN(n90) );
  NAND4_X1 U51 ( .A1(n62), .A2(n177), .A3(n57), .A4(n180), .ZN(n65) );
  NAND2_X1 U52 ( .A1(n169), .A2(n63), .ZN(n60) );
  NAND3_X1 U53 ( .A1(s_tick), .A2(n64), .A3(U27_DATA2_0), .ZN(n63) );
  INV_X1 U54 ( .A(n67), .ZN(n169) );
  OAI21_X1 U55 ( .B1(rx), .B2(n39), .A(n68), .ZN(n67) );
  INV_X1 U56 ( .A(n32), .ZN(n171) );
  AOI22_X1 U57 ( .A1(n33), .A2(U22_DATA1_0), .B1(n173), .B2(n34), .ZN(n32) );
  OAI21_X1 U58 ( .B1(n37), .B2(n38), .A(n36), .ZN(n33) );
  AND2_X1 U59 ( .A1(n35), .A2(n36), .ZN(n34) );
  OAI22_X1 U60 ( .A1(n41), .A2(n7), .B1(n170), .B2(n6), .ZN(n81) );
  OAI22_X1 U61 ( .A1(n41), .A2(n6), .B1(n170), .B2(n5), .ZN(n80) );
  OAI22_X1 U62 ( .A1(n41), .A2(n5), .B1(n170), .B2(n4), .ZN(n79) );
  OAI22_X1 U63 ( .A1(n41), .A2(n4), .B1(n170), .B2(n3), .ZN(n78) );
  OAI22_X1 U64 ( .A1(n41), .A2(n3), .B1(n170), .B2(n2), .ZN(n77) );
  OAI22_X1 U65 ( .A1(n41), .A2(n2), .B1(n170), .B2(n1), .ZN(n76) );
  OAI21_X1 U66 ( .B1(n170), .B2(n7), .A(n42), .ZN(n82) );
  NAND2_X1 U67 ( .A1(data_out[0]), .A2(n170), .ZN(n42) );
  AND4_X1 U68 ( .A1(n166), .A2(n30), .A3(n29), .A4(n28), .ZN(n56) );
  NAND4_X1 U69 ( .A1(U3_U3_DATA3_3), .A2(U3_U3_DATA3_2), .A3(U3_U3_DATA3_1), 
        .A4(U3_U3_DATA3_0), .ZN(n64) );
  NAND2_X1 U70 ( .A1(U27_DATA2_1), .A2(n18), .ZN(n37) );
  NAND2_X1 U71 ( .A1(U27_DATA2_0), .A2(U27_DATA2_1), .ZN(n69) );
  OAI22_X1 U72 ( .A1(n73), .A2(n30), .B1(n74), .B2(n26), .ZN(n48) );
  OAI22_X1 U73 ( .A1(n73), .A2(n29), .B1(n74), .B2(n25), .ZN(n50) );
  AOI22_X1 U74 ( .A1(n173), .A2(U3_U3_DATA4_2), .B1(n174), .B2(U3_U3_DATA3_2), 
        .ZN(n52) );
  INV_X1 U75 ( .A(n74), .ZN(n174) );
  XNOR2_X1 U76 ( .A(n71), .B(n72), .ZN(n58) );
  OAI22_X1 U77 ( .A1(n27), .A2(n73), .B1(n74), .B2(n19), .ZN(n71) );
  NOR2_X1 U78 ( .A1(n52), .A2(n51), .ZN(n72) );
  NAND2_X1 U79 ( .A1(U27_DATA2_0), .A2(n13), .ZN(n70) );
endmodule


module dual_gray_counter_addr_size8_2_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[8]), .B(A[8]), .Z(SUM[8]) );
endmodule


module dual_gray_counter_addr_size8_2 ( clk, gray_count_st, gray_count_nd, 
        reset_n, en );
  output [8:0] gray_count_st;
  output [7:0] gray_count_nd;
  input clk, reset_n, en;
  wire   n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54;
  wire   [7:0] Q_reg;
  wire   [8:0] Q_next;
  assign gray_count_nd[6] = gray_count_st[6];
  assign gray_count_nd[5] = gray_count_st[5];
  assign gray_count_nd[4] = gray_count_st[4];
  assign gray_count_nd[3] = gray_count_st[3];
  assign gray_count_nd[2] = gray_count_st[2];
  assign gray_count_nd[1] = gray_count_st[1];
  assign gray_count_nd[0] = gray_count_st[0];

  DFFR_X1 Q_reg_reg_0_ ( .D(n28), .CK(clk), .RN(reset_n), .Q(Q_reg[0]), .QN(
        n37) );
  DFFR_X1 Q_reg_reg_1_ ( .D(n29), .CK(clk), .RN(reset_n), .Q(Q_reg[1]), .QN(
        n38) );
  DFFR_X1 Q_reg_reg_2_ ( .D(n30), .CK(clk), .RN(reset_n), .Q(Q_reg[2]), .QN(
        n39) );
  DFFR_X1 Q_reg_reg_3_ ( .D(n31), .CK(clk), .RN(reset_n), .Q(Q_reg[3]), .QN(
        n40) );
  DFFR_X1 Q_reg_reg_4_ ( .D(n32), .CK(clk), .RN(reset_n), .Q(Q_reg[4]), .QN(
        n41) );
  DFFR_X1 Q_reg_reg_5_ ( .D(n33), .CK(clk), .RN(reset_n), .Q(Q_reg[5]), .QN(
        n42) );
  DFFR_X1 Q_reg_reg_6_ ( .D(n34), .CK(clk), .RN(reset_n), .Q(Q_reg[6]), .QN(
        n43) );
  DFFR_X1 Q_reg_reg_7_ ( .D(n35), .CK(clk), .RN(reset_n), .Q(Q_reg[7]), .QN(
        n44) );
  DFFR_X1 Q_reg_reg_8_ ( .D(n36), .CK(clk), .RN(reset_n), .Q(gray_count_st[8]), 
        .QN(n45) );
  XOR2_X1 U21 ( .A(n44), .B(n43), .Z(gray_count_st[6]) );
  XOR2_X1 U22 ( .A(n43), .B(n42), .Z(gray_count_st[5]) );
  XOR2_X1 U23 ( .A(n42), .B(n41), .Z(gray_count_st[4]) );
  XOR2_X1 U24 ( .A(n41), .B(n40), .Z(gray_count_st[3]) );
  XOR2_X1 U25 ( .A(n40), .B(n39), .Z(gray_count_st[2]) );
  XOR2_X1 U26 ( .A(n39), .B(n38), .Z(gray_count_st[1]) );
  XOR2_X1 U27 ( .A(n38), .B(n37), .Z(gray_count_st[0]) );
  XOR2_X1 U29 ( .A(n44), .B(n45), .Z(gray_count_st[7]) );
  dual_gray_counter_addr_size8_2_DW01_inc_0 add_48 ( .A({gray_count_st[8], 
        Q_reg}), .SUM(Q_next) );
  XNOR2_X1 U3 ( .A(n45), .B(gray_count_st[7]), .ZN(gray_count_nd[7]) );
  OAI21_X1 U4 ( .B1(n45), .B2(en), .A(n54), .ZN(n36) );
  NAND2_X1 U5 ( .A1(en), .A2(Q_next[8]), .ZN(n54) );
  OAI21_X1 U6 ( .B1(n44), .B2(en), .A(n53), .ZN(n35) );
  NAND2_X1 U7 ( .A1(Q_next[7]), .A2(en), .ZN(n53) );
  OAI21_X1 U8 ( .B1(n43), .B2(en), .A(n52), .ZN(n34) );
  NAND2_X1 U9 ( .A1(Q_next[6]), .A2(en), .ZN(n52) );
  OAI21_X1 U10 ( .B1(n42), .B2(en), .A(n51), .ZN(n33) );
  NAND2_X1 U11 ( .A1(Q_next[5]), .A2(en), .ZN(n51) );
  OAI21_X1 U12 ( .B1(n41), .B2(en), .A(n50), .ZN(n32) );
  NAND2_X1 U13 ( .A1(Q_next[4]), .A2(en), .ZN(n50) );
  OAI21_X1 U14 ( .B1(n40), .B2(en), .A(n49), .ZN(n31) );
  NAND2_X1 U15 ( .A1(Q_next[3]), .A2(en), .ZN(n49) );
  OAI21_X1 U16 ( .B1(n39), .B2(en), .A(n48), .ZN(n30) );
  NAND2_X1 U17 ( .A1(Q_next[2]), .A2(en), .ZN(n48) );
  OAI21_X1 U18 ( .B1(n38), .B2(en), .A(n47), .ZN(n29) );
  NAND2_X1 U19 ( .A1(Q_next[1]), .A2(en), .ZN(n47) );
  OAI21_X1 U20 ( .B1(n37), .B2(en), .A(n46), .ZN(n28) );
  NAND2_X1 U28 ( .A1(Q_next[0]), .A2(en), .ZN(n46) );
endmodule


module dual_gray_counter_addr_size8_0 ( clk, gray_count_st, gray_count_nd, 
        reset_n, en );
  output [8:0] gray_count_st;
  output [7:0] gray_count_nd;
  input clk, reset_n, en;
  wire   n2, n3, n4, n6, n7, n9, n10, n12, n14, n15, n17, n19, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n1, n5, n8, n11;
  assign gray_count_nd[6] = gray_count_st[6];
  assign gray_count_nd[5] = gray_count_st[5];
  assign gray_count_nd[4] = gray_count_st[4];
  assign gray_count_nd[3] = gray_count_st[3];
  assign gray_count_nd[2] = gray_count_st[2];
  assign gray_count_nd[1] = gray_count_st[1];
  assign gray_count_nd[0] = gray_count_st[0];

  XOR2_X1 U3 ( .A(gray_count_st[8]), .B(n2), .Z(n22) );
  XOR2_X1 U5 ( .A(n3), .B(n15), .Z(n23) );
  XOR2_X1 U7 ( .A(n4), .B(n11), .Z(n24) );
  XOR2_X1 U9 ( .A(n6), .B(n17), .Z(n25) );
  XOR2_X1 U11 ( .A(n7), .B(n8), .Z(n26) );
  XOR2_X1 U13 ( .A(n9), .B(n19), .Z(n27) );
  XOR2_X1 U15 ( .A(n10), .B(n5), .Z(n28) );
  XOR2_X1 U17 ( .A(n12), .B(n21), .Z(n29) );
  XOR2_X1 U19 ( .A(en), .B(n1), .Z(n30) );
  XOR2_X1 U31 ( .A(gray_count_st[8]), .B(gray_count_st[7]), .Z(
        gray_count_nd[7]) );
  XOR2_X1 U32 ( .A(n14), .B(n15), .Z(gray_count_st[7]) );
  DFFR_X1 Q_reg_reg_0_ ( .D(n30), .CK(clk), .RN(reset_n), .Q(n1) );
  DFFR_X1 Q_reg_reg_1_ ( .D(n29), .CK(clk), .RN(reset_n), .QN(n21) );
  DFFR_X1 Q_reg_reg_2_ ( .D(n28), .CK(clk), .RN(reset_n), .Q(n5) );
  DFFR_X1 Q_reg_reg_3_ ( .D(n27), .CK(clk), .RN(reset_n), .QN(n19) );
  DFFR_X1 Q_reg_reg_4_ ( .D(n26), .CK(clk), .RN(reset_n), .Q(n8) );
  DFFR_X1 Q_reg_reg_5_ ( .D(n25), .CK(clk), .RN(reset_n), .QN(n17) );
  DFFR_X1 Q_reg_reg_6_ ( .D(n24), .CK(clk), .RN(reset_n), .Q(n11) );
  DFFR_X1 Q_reg_reg_7_ ( .D(n23), .CK(clk), .RN(reset_n), .QN(n15) );
  DFFR_X1 Q_reg_reg_8_ ( .D(n22), .CK(clk), .RN(reset_n), .Q(gray_count_st[8]), 
        .QN(n14) );
  NAND2_X1 U4 ( .A1(en), .A2(n1), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n4), .A2(n11), .ZN(n3) );
  NAND2_X1 U8 ( .A1(n10), .A2(n5), .ZN(n9) );
  NAND2_X1 U10 ( .A1(n7), .A2(n8), .ZN(n6) );
  NOR2_X1 U12 ( .A1(n12), .A2(n21), .ZN(n10) );
  NOR2_X1 U14 ( .A1(n9), .A2(n19), .ZN(n7) );
  NOR2_X1 U16 ( .A1(n6), .A2(n17), .ZN(n4) );
  NOR2_X1 U18 ( .A1(n15), .A2(n3), .ZN(n2) );
  XNOR2_X1 U20 ( .A(n11), .B(n17), .ZN(gray_count_st[5]) );
  XNOR2_X1 U21 ( .A(n17), .B(n8), .ZN(gray_count_st[4]) );
  XNOR2_X1 U22 ( .A(n8), .B(n19), .ZN(gray_count_st[3]) );
  XNOR2_X1 U23 ( .A(n5), .B(n21), .ZN(gray_count_st[1]) );
  XNOR2_X1 U24 ( .A(n19), .B(n5), .ZN(gray_count_st[2]) );
  XNOR2_X1 U25 ( .A(n21), .B(n1), .ZN(gray_count_st[0]) );
  XNOR2_X1 U26 ( .A(n15), .B(n11), .ZN(gray_count_st[6]) );
endmodule


module fifo_control_unit_addr_size8_0 ( reset_n, w_clk, r_clk, rd, wr, addr_r, 
        addr_w, full, empty, we_enable, rd_enable );
  output [7:0] addr_r;
  output [7:0] addr_w;
  input reset_n, w_clk, r_clk, rd, wr;
  output full, empty, we_enable, rd_enable;
  wire   eq_127_B_0_, eq_127_B_1_, eq_127_B_2_, eq_127_B_3_, eq_127_B_4_,
         eq_127_B_5_, eq_127_B_6_, eq_127_B_7_, eq_127_B_8_, eq_127_A_0_,
         eq_127_A_1_, eq_127_A_2_, eq_127_A_3_, eq_127_A_4_, eq_127_A_5_,
         eq_127_A_6_, eq_127_A_7_, eq_127_A_8_, eq_117_B_0_, eq_117_B_1_,
         eq_117_B_2_, eq_117_B_3_, eq_117_B_4_, eq_117_B_5_, eq_117_B_6_,
         eq_117_A_0_, eq_117_A_1_, eq_117_A_2_, eq_117_A_3_, eq_117_A_4_,
         eq_117_A_5_, eq_117_A_6_, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [8:7] ptr_w;
  wire   [8:0] ptr_w_syn_1;
  wire   [8:7] ptr_r_syn;
  wire   [8:0] ptr_r_syn_1;

  XOR2_X1 U19 ( .A(eq_117_B_6_), .B(eq_117_A_6_), .Z(n12) );
  XOR2_X1 U20 ( .A(eq_117_B_2_), .B(eq_117_A_2_), .Z(n11) );
  XOR2_X1 U21 ( .A(eq_117_B_1_), .B(eq_117_A_1_), .Z(n10) );
  XOR2_X1 U22 ( .A(eq_117_B_0_), .B(eq_117_A_0_), .Z(n9) );
  XOR2_X1 U23 ( .A(eq_117_B_3_), .B(eq_117_A_3_), .Z(n13) );
  XOR2_X1 U24 ( .A(eq_127_B_8_), .B(eq_127_A_8_), .Z(n23) );
  XOR2_X1 U25 ( .A(eq_127_B_7_), .B(eq_127_A_7_), .Z(n22) );
  XOR2_X1 U26 ( .A(eq_127_B_6_), .B(eq_127_A_6_), .Z(n21) );
  XOR2_X1 U27 ( .A(eq_127_B_5_), .B(eq_127_A_5_), .Z(n20) );
  XOR2_X1 U28 ( .A(eq_127_B_1_), .B(eq_127_A_1_), .Z(n26) );
  XOR2_X1 U29 ( .A(eq_127_B_0_), .B(eq_127_A_0_), .Z(n25) );
  XOR2_X1 U30 ( .A(eq_127_B_2_), .B(eq_127_A_2_), .Z(n24) );
  dual_gray_counter_addr_size8_2 read_ptr ( .clk(r_clk), .gray_count_st({
        eq_127_B_8_, eq_127_B_7_, eq_127_B_6_, eq_127_B_5_, eq_127_B_4_, 
        eq_127_B_3_, eq_127_B_2_, eq_127_B_1_, eq_127_B_0_}), .gray_count_nd(
        addr_r), .reset_n(reset_n), .en(rd_enable) );
  dual_gray_counter_addr_size8_0 write_ptr ( .clk(w_clk), .gray_count_st({
        ptr_w, eq_117_A_6_, eq_117_A_5_, eq_117_A_4_, eq_117_A_3_, eq_117_A_2_, 
        eq_117_A_1_, eq_117_A_0_}), .gray_count_nd(addr_w), .reset_n(reset_n), 
        .en(we_enable) );
  DFFR_X1 ptr_w_syn_reg_8_ ( .D(ptr_w_syn_1[8]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_8_) );
  DFFR_X1 ptr_w_syn_reg_7_ ( .D(ptr_w_syn_1[7]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_7_) );
  DFFR_X1 ptr_w_syn_reg_6_ ( .D(ptr_w_syn_1[6]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_6_) );
  DFFR_X1 ptr_w_syn_reg_5_ ( .D(ptr_w_syn_1[5]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_5_) );
  DFFR_X1 ptr_w_syn_reg_4_ ( .D(ptr_w_syn_1[4]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_4_) );
  DFFR_X1 ptr_w_syn_reg_3_ ( .D(ptr_w_syn_1[3]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_3_) );
  DFFR_X1 ptr_w_syn_reg_2_ ( .D(ptr_w_syn_1[2]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_2_) );
  DFFR_X1 ptr_w_syn_reg_1_ ( .D(ptr_w_syn_1[1]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_1_) );
  DFFR_X1 ptr_w_syn_reg_0_ ( .D(ptr_w_syn_1[0]), .CK(r_clk), .RN(reset_n), .Q(
        eq_127_A_0_) );
  DFFR_X1 ptr_r_syn_reg_8_ ( .D(ptr_r_syn_1[8]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[8]) );
  DFFR_X1 ptr_r_syn_reg_7_ ( .D(ptr_r_syn_1[7]), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn[7]) );
  DFFR_X1 ptr_r_syn_reg_6_ ( .D(ptr_r_syn_1[6]), .CK(w_clk), .RN(reset_n), .Q(
        eq_117_B_6_) );
  DFFR_X1 ptr_r_syn_reg_5_ ( .D(ptr_r_syn_1[5]), .CK(w_clk), .RN(reset_n), .Q(
        eq_117_B_5_) );
  DFFR_X1 ptr_r_syn_reg_4_ ( .D(ptr_r_syn_1[4]), .CK(w_clk), .RN(reset_n), .Q(
        eq_117_B_4_) );
  DFFR_X1 ptr_r_syn_reg_3_ ( .D(ptr_r_syn_1[3]), .CK(w_clk), .RN(reset_n), .Q(
        eq_117_B_3_) );
  DFFR_X1 ptr_r_syn_reg_2_ ( .D(ptr_r_syn_1[2]), .CK(w_clk), .RN(reset_n), .Q(
        eq_117_B_2_) );
  DFFR_X1 ptr_r_syn_reg_1_ ( .D(ptr_r_syn_1[1]), .CK(w_clk), .RN(reset_n), .Q(
        eq_117_B_1_) );
  DFFR_X1 ptr_r_syn_reg_0_ ( .D(ptr_r_syn_1[0]), .CK(w_clk), .RN(reset_n), .Q(
        eq_117_B_0_) );
  DFFR_X1 ptr_w_syn_1_reg_8_ ( .D(ptr_w[8]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[8]) );
  DFFR_X1 ptr_r_syn_1_reg_8_ ( .D(eq_127_B_8_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[8]) );
  DFFR_X1 ptr_r_syn_1_reg_7_ ( .D(eq_127_B_7_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[7]) );
  DFFR_X1 ptr_w_syn_1_reg_7_ ( .D(ptr_w[7]), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[7]) );
  DFFR_X1 ptr_r_syn_1_reg_4_ ( .D(eq_127_B_4_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[4]) );
  DFFR_X1 ptr_w_syn_1_reg_0_ ( .D(eq_117_A_0_), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[0]) );
  DFFR_X1 ptr_r_syn_1_reg_5_ ( .D(eq_127_B_5_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[5]) );
  DFFR_X1 ptr_r_syn_1_reg_6_ ( .D(eq_127_B_6_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[6]) );
  DFFR_X1 ptr_w_syn_1_reg_3_ ( .D(eq_117_A_3_), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[3]) );
  DFFR_X1 ptr_w_syn_1_reg_1_ ( .D(eq_117_A_1_), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[1]) );
  DFFR_X1 ptr_w_syn_1_reg_4_ ( .D(eq_117_A_4_), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[4]) );
  DFFR_X1 ptr_w_syn_1_reg_5_ ( .D(eq_117_A_5_), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[5]) );
  DFFR_X1 ptr_r_syn_1_reg_3_ ( .D(eq_127_B_3_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[3]) );
  DFFR_X1 ptr_r_syn_1_reg_2_ ( .D(eq_127_B_2_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[2]) );
  DFFR_X1 ptr_w_syn_1_reg_6_ ( .D(eq_117_A_6_), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[6]) );
  DFFR_X1 ptr_w_syn_1_reg_2_ ( .D(eq_117_A_2_), .CK(r_clk), .RN(reset_n), .Q(
        ptr_w_syn_1[2]) );
  DFFR_X1 ptr_r_syn_1_reg_0_ ( .D(eq_127_B_0_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[0]) );
  DFFR_X1 ptr_r_syn_1_reg_1_ ( .D(eq_127_B_1_), .CK(w_clk), .RN(reset_n), .Q(
        ptr_r_syn_1[1]) );
  AND2_X1 U3 ( .A1(wr), .A2(n3), .ZN(we_enable) );
  INV_X1 U4 ( .A(n4), .ZN(empty) );
  INV_X1 U5 ( .A(n3), .ZN(full) );
  AND2_X1 U6 ( .A1(rd), .A2(n4), .ZN(rd_enable) );
  NOR3_X1 U7 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n18) );
  NAND4_X1 U8 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n4) );
  XNOR2_X1 U9 ( .A(eq_127_B_4_), .B(eq_127_A_4_), .ZN(n16) );
  XNOR2_X1 U10 ( .A(eq_127_B_3_), .B(eq_127_A_3_), .ZN(n17) );
  NOR4_X1 U11 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  NOR4_X1 U12 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n8) );
  NAND4_X1 U13 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n3) );
  XNOR2_X1 U14 ( .A(eq_117_B_5_), .B(eq_117_A_5_), .ZN(n5) );
  XNOR2_X1 U15 ( .A(eq_117_B_4_), .B(eq_117_A_4_), .ZN(n6) );
  NOR3_X1 U16 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n7) );
  XNOR2_X1 U17 ( .A(ptr_w[7]), .B(ptr_r_syn[7]), .ZN(n15) );
  XNOR2_X1 U18 ( .A(ptr_w[8]), .B(ptr_r_syn[8]), .ZN(n14) );
endmodule


module reg_memory_file_addr_size8_word_width8_0 ( we_s, clk, addr_r, addr_w, 
        data_w, data_r );
  input [7:0] addr_r;
  input [7:0] addr_w;
  input [7:0] data_w;
  output [7:0] data_r;
  input we_s, clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258;
  wire   [2608:577] n;

  DFF_X1 reg_mem_reg_0__7_ ( .D(n7103), .CK(clk), .Q(n[2608]), .QN(n1) );
  DFF_X1 reg_mem_reg_0__6_ ( .D(n7102), .CK(clk), .Q(n[2607]), .QN(n2) );
  DFF_X1 reg_mem_reg_0__5_ ( .D(n7101), .CK(clk), .Q(n[2606]), .QN(n3) );
  DFF_X1 reg_mem_reg_0__4_ ( .D(n7100), .CK(clk), .Q(n[2605]), .QN(n4) );
  DFF_X1 reg_mem_reg_0__3_ ( .D(n7099), .CK(clk), .Q(n[2604]), .QN(n5) );
  DFF_X1 reg_mem_reg_0__2_ ( .D(n7098), .CK(clk), .Q(n[2603]), .QN(n6) );
  DFF_X1 reg_mem_reg_0__1_ ( .D(n7097), .CK(clk), .Q(n[2602]), .QN(n7) );
  DFF_X1 reg_mem_reg_0__0_ ( .D(n7096), .CK(clk), .Q(n[2601]), .QN(n8) );
  DFF_X1 reg_mem_reg_1__7_ ( .D(n7095), .CK(clk), .Q(n[2600]), .QN(n9) );
  DFF_X1 reg_mem_reg_1__6_ ( .D(n7094), .CK(clk), .Q(n[2599]), .QN(n10) );
  DFF_X1 reg_mem_reg_1__5_ ( .D(n7093), .CK(clk), .Q(n[2598]), .QN(n11) );
  DFF_X1 reg_mem_reg_1__4_ ( .D(n7092), .CK(clk), .Q(n[2597]), .QN(n12) );
  DFF_X1 reg_mem_reg_1__3_ ( .D(n7091), .CK(clk), .Q(n[2596]), .QN(n13) );
  DFF_X1 reg_mem_reg_1__2_ ( .D(n7090), .CK(clk), .Q(n[2595]), .QN(n14) );
  DFF_X1 reg_mem_reg_1__1_ ( .D(n7089), .CK(clk), .Q(n[2594]), .QN(n15) );
  DFF_X1 reg_mem_reg_1__0_ ( .D(n7088), .CK(clk), .Q(n[2593]), .QN(n16) );
  DFF_X1 reg_mem_reg_2__7_ ( .D(n7087), .CK(clk), .QN(n17) );
  DFF_X1 reg_mem_reg_2__6_ ( .D(n7086), .CK(clk), .QN(n18) );
  DFF_X1 reg_mem_reg_2__5_ ( .D(n7085), .CK(clk), .QN(n19) );
  DFF_X1 reg_mem_reg_2__4_ ( .D(n7084), .CK(clk), .QN(n20) );
  DFF_X1 reg_mem_reg_2__3_ ( .D(n7083), .CK(clk), .QN(n21) );
  DFF_X1 reg_mem_reg_2__2_ ( .D(n7082), .CK(clk), .QN(n22) );
  DFF_X1 reg_mem_reg_2__1_ ( .D(n7081), .CK(clk), .QN(n23) );
  DFF_X1 reg_mem_reg_2__0_ ( .D(n7080), .CK(clk), .QN(n24) );
  DFF_X1 reg_mem_reg_3__7_ ( .D(n7079), .CK(clk), .QN(n25) );
  DFF_X1 reg_mem_reg_3__6_ ( .D(n7078), .CK(clk), .QN(n26) );
  DFF_X1 reg_mem_reg_3__5_ ( .D(n7077), .CK(clk), .QN(n27) );
  DFF_X1 reg_mem_reg_3__4_ ( .D(n7076), .CK(clk), .QN(n28) );
  DFF_X1 reg_mem_reg_3__3_ ( .D(n7075), .CK(clk), .QN(n29) );
  DFF_X1 reg_mem_reg_3__2_ ( .D(n7074), .CK(clk), .QN(n30) );
  DFF_X1 reg_mem_reg_3__1_ ( .D(n7073), .CK(clk), .QN(n31) );
  DFF_X1 reg_mem_reg_3__0_ ( .D(n7072), .CK(clk), .QN(n32) );
  DFF_X1 reg_mem_reg_4__7_ ( .D(n7071), .CK(clk), .Q(n[2576]), .QN(n33) );
  DFF_X1 reg_mem_reg_4__6_ ( .D(n7070), .CK(clk), .Q(n[2575]), .QN(n34) );
  DFF_X1 reg_mem_reg_4__5_ ( .D(n7069), .CK(clk), .Q(n[2574]), .QN(n35) );
  DFF_X1 reg_mem_reg_4__4_ ( .D(n7068), .CK(clk), .Q(n[2573]), .QN(n36) );
  DFF_X1 reg_mem_reg_4__3_ ( .D(n7067), .CK(clk), .Q(n[2572]), .QN(n37) );
  DFF_X1 reg_mem_reg_4__2_ ( .D(n7066), .CK(clk), .Q(n[2571]), .QN(n38) );
  DFF_X1 reg_mem_reg_4__1_ ( .D(n7065), .CK(clk), .Q(n[2570]), .QN(n39) );
  DFF_X1 reg_mem_reg_4__0_ ( .D(n7064), .CK(clk), .Q(n[2569]), .QN(n40) );
  DFF_X1 reg_mem_reg_5__7_ ( .D(n7063), .CK(clk), .Q(n[2568]), .QN(n41) );
  DFF_X1 reg_mem_reg_5__6_ ( .D(n7062), .CK(clk), .Q(n[2567]), .QN(n42) );
  DFF_X1 reg_mem_reg_5__5_ ( .D(n7061), .CK(clk), .Q(n[2566]), .QN(n43) );
  DFF_X1 reg_mem_reg_5__4_ ( .D(n7060), .CK(clk), .Q(n[2565]), .QN(n44) );
  DFF_X1 reg_mem_reg_5__3_ ( .D(n7059), .CK(clk), .Q(n[2564]), .QN(n45) );
  DFF_X1 reg_mem_reg_5__2_ ( .D(n7058), .CK(clk), .Q(n[2563]), .QN(n46) );
  DFF_X1 reg_mem_reg_5__1_ ( .D(n7057), .CK(clk), .Q(n[2562]), .QN(n47) );
  DFF_X1 reg_mem_reg_5__0_ ( .D(n7056), .CK(clk), .Q(n[2561]), .QN(n48) );
  DFF_X1 reg_mem_reg_6__7_ ( .D(n7055), .CK(clk), .QN(n49) );
  DFF_X1 reg_mem_reg_6__6_ ( .D(n7054), .CK(clk), .QN(n50) );
  DFF_X1 reg_mem_reg_6__5_ ( .D(n7053), .CK(clk), .QN(n51) );
  DFF_X1 reg_mem_reg_6__4_ ( .D(n7052), .CK(clk), .QN(n52) );
  DFF_X1 reg_mem_reg_6__3_ ( .D(n7051), .CK(clk), .QN(n53) );
  DFF_X1 reg_mem_reg_6__2_ ( .D(n7050), .CK(clk), .QN(n54) );
  DFF_X1 reg_mem_reg_6__1_ ( .D(n7049), .CK(clk), .QN(n55) );
  DFF_X1 reg_mem_reg_6__0_ ( .D(n7048), .CK(clk), .QN(n56) );
  DFF_X1 reg_mem_reg_7__7_ ( .D(n7047), .CK(clk), .QN(n57) );
  DFF_X1 reg_mem_reg_7__6_ ( .D(n7046), .CK(clk), .QN(n58) );
  DFF_X1 reg_mem_reg_7__5_ ( .D(n7045), .CK(clk), .QN(n59) );
  DFF_X1 reg_mem_reg_7__4_ ( .D(n7044), .CK(clk), .QN(n60) );
  DFF_X1 reg_mem_reg_7__3_ ( .D(n7043), .CK(clk), .QN(n61) );
  DFF_X1 reg_mem_reg_7__2_ ( .D(n7042), .CK(clk), .QN(n62) );
  DFF_X1 reg_mem_reg_7__1_ ( .D(n7041), .CK(clk), .QN(n63) );
  DFF_X1 reg_mem_reg_7__0_ ( .D(n7040), .CK(clk), .QN(n64) );
  DFF_X1 reg_mem_reg_8__7_ ( .D(n7039), .CK(clk), .Q(n[2544]), .QN(n65) );
  DFF_X1 reg_mem_reg_8__6_ ( .D(n7038), .CK(clk), .Q(n[2543]), .QN(n66) );
  DFF_X1 reg_mem_reg_8__5_ ( .D(n7037), .CK(clk), .Q(n[2542]), .QN(n67) );
  DFF_X1 reg_mem_reg_8__4_ ( .D(n7036), .CK(clk), .Q(n[2541]), .QN(n68) );
  DFF_X1 reg_mem_reg_8__3_ ( .D(n7035), .CK(clk), .Q(n[2540]), .QN(n69) );
  DFF_X1 reg_mem_reg_8__2_ ( .D(n7034), .CK(clk), .Q(n[2539]), .QN(n70) );
  DFF_X1 reg_mem_reg_8__1_ ( .D(n7033), .CK(clk), .Q(n[2538]), .QN(n71) );
  DFF_X1 reg_mem_reg_8__0_ ( .D(n7032), .CK(clk), .Q(n[2537]), .QN(n72) );
  DFF_X1 reg_mem_reg_9__7_ ( .D(n7031), .CK(clk), .Q(n[2536]), .QN(n73) );
  DFF_X1 reg_mem_reg_9__6_ ( .D(n7030), .CK(clk), .Q(n[2535]), .QN(n74) );
  DFF_X1 reg_mem_reg_9__5_ ( .D(n7029), .CK(clk), .Q(n[2534]), .QN(n75) );
  DFF_X1 reg_mem_reg_9__4_ ( .D(n7028), .CK(clk), .Q(n[2533]), .QN(n76) );
  DFF_X1 reg_mem_reg_9__3_ ( .D(n7027), .CK(clk), .Q(n[2532]), .QN(n77) );
  DFF_X1 reg_mem_reg_9__2_ ( .D(n7026), .CK(clk), .Q(n[2531]), .QN(n78) );
  DFF_X1 reg_mem_reg_9__1_ ( .D(n7025), .CK(clk), .Q(n[2530]), .QN(n79) );
  DFF_X1 reg_mem_reg_9__0_ ( .D(n7024), .CK(clk), .Q(n[2529]), .QN(n80) );
  DFF_X1 reg_mem_reg_10__7_ ( .D(n7023), .CK(clk), .QN(n81) );
  DFF_X1 reg_mem_reg_10__6_ ( .D(n7022), .CK(clk), .QN(n82) );
  DFF_X1 reg_mem_reg_10__5_ ( .D(n7021), .CK(clk), .QN(n83) );
  DFF_X1 reg_mem_reg_10__4_ ( .D(n7020), .CK(clk), .QN(n84) );
  DFF_X1 reg_mem_reg_10__3_ ( .D(n7019), .CK(clk), .QN(n85) );
  DFF_X1 reg_mem_reg_10__2_ ( .D(n7018), .CK(clk), .QN(n86) );
  DFF_X1 reg_mem_reg_10__1_ ( .D(n7017), .CK(clk), .QN(n87) );
  DFF_X1 reg_mem_reg_10__0_ ( .D(n7016), .CK(clk), .QN(n88) );
  DFF_X1 reg_mem_reg_11__7_ ( .D(n7015), .CK(clk), .QN(n89) );
  DFF_X1 reg_mem_reg_11__6_ ( .D(n7014), .CK(clk), .QN(n90) );
  DFF_X1 reg_mem_reg_11__5_ ( .D(n7013), .CK(clk), .QN(n91) );
  DFF_X1 reg_mem_reg_11__4_ ( .D(n7012), .CK(clk), .QN(n92) );
  DFF_X1 reg_mem_reg_11__3_ ( .D(n7011), .CK(clk), .QN(n93) );
  DFF_X1 reg_mem_reg_11__2_ ( .D(n7010), .CK(clk), .QN(n94) );
  DFF_X1 reg_mem_reg_11__1_ ( .D(n7009), .CK(clk), .QN(n95) );
  DFF_X1 reg_mem_reg_11__0_ ( .D(n7008), .CK(clk), .QN(n96) );
  DFF_X1 reg_mem_reg_12__7_ ( .D(n7007), .CK(clk), .Q(n[2512]), .QN(n97) );
  DFF_X1 reg_mem_reg_12__6_ ( .D(n7006), .CK(clk), .Q(n[2511]), .QN(n98) );
  DFF_X1 reg_mem_reg_12__5_ ( .D(n7005), .CK(clk), .Q(n[2510]), .QN(n99) );
  DFF_X1 reg_mem_reg_12__4_ ( .D(n7004), .CK(clk), .Q(n[2509]), .QN(n100) );
  DFF_X1 reg_mem_reg_12__3_ ( .D(n7003), .CK(clk), .Q(n[2508]), .QN(n101) );
  DFF_X1 reg_mem_reg_12__2_ ( .D(n7002), .CK(clk), .Q(n[2507]), .QN(n102) );
  DFF_X1 reg_mem_reg_12__1_ ( .D(n7001), .CK(clk), .Q(n[2506]), .QN(n103) );
  DFF_X1 reg_mem_reg_12__0_ ( .D(n7000), .CK(clk), .Q(n[2505]), .QN(n104) );
  DFF_X1 reg_mem_reg_13__7_ ( .D(n6999), .CK(clk), .Q(n[2504]), .QN(n105) );
  DFF_X1 reg_mem_reg_13__6_ ( .D(n6998), .CK(clk), .Q(n[2503]), .QN(n106) );
  DFF_X1 reg_mem_reg_13__5_ ( .D(n6997), .CK(clk), .Q(n[2502]), .QN(n107) );
  DFF_X1 reg_mem_reg_13__4_ ( .D(n6996), .CK(clk), .Q(n[2501]), .QN(n108) );
  DFF_X1 reg_mem_reg_13__3_ ( .D(n6995), .CK(clk), .Q(n[2500]), .QN(n109) );
  DFF_X1 reg_mem_reg_13__2_ ( .D(n6994), .CK(clk), .Q(n[2499]), .QN(n110) );
  DFF_X1 reg_mem_reg_13__1_ ( .D(n6993), .CK(clk), .Q(n[2498]), .QN(n111) );
  DFF_X1 reg_mem_reg_13__0_ ( .D(n6992), .CK(clk), .Q(n[2497]), .QN(n112) );
  DFF_X1 reg_mem_reg_14__7_ ( .D(n6991), .CK(clk), .QN(n113) );
  DFF_X1 reg_mem_reg_14__6_ ( .D(n6990), .CK(clk), .QN(n114) );
  DFF_X1 reg_mem_reg_14__5_ ( .D(n6989), .CK(clk), .QN(n115) );
  DFF_X1 reg_mem_reg_14__4_ ( .D(n6988), .CK(clk), .QN(n116) );
  DFF_X1 reg_mem_reg_14__3_ ( .D(n6987), .CK(clk), .QN(n117) );
  DFF_X1 reg_mem_reg_14__2_ ( .D(n6986), .CK(clk), .QN(n118) );
  DFF_X1 reg_mem_reg_14__1_ ( .D(n6985), .CK(clk), .QN(n119) );
  DFF_X1 reg_mem_reg_14__0_ ( .D(n6984), .CK(clk), .QN(n120) );
  DFF_X1 reg_mem_reg_15__7_ ( .D(n6983), .CK(clk), .QN(n121) );
  DFF_X1 reg_mem_reg_15__6_ ( .D(n6982), .CK(clk), .QN(n122) );
  DFF_X1 reg_mem_reg_15__5_ ( .D(n6981), .CK(clk), .QN(n123) );
  DFF_X1 reg_mem_reg_15__4_ ( .D(n6980), .CK(clk), .QN(n124) );
  DFF_X1 reg_mem_reg_15__3_ ( .D(n6979), .CK(clk), .QN(n125) );
  DFF_X1 reg_mem_reg_15__2_ ( .D(n6978), .CK(clk), .QN(n126) );
  DFF_X1 reg_mem_reg_15__1_ ( .D(n6977), .CK(clk), .QN(n127) );
  DFF_X1 reg_mem_reg_15__0_ ( .D(n6976), .CK(clk), .QN(n128) );
  DFF_X1 reg_mem_reg_16__7_ ( .D(n6975), .CK(clk), .Q(n[2480]), .QN(n129) );
  DFF_X1 reg_mem_reg_16__6_ ( .D(n6974), .CK(clk), .Q(n[2479]), .QN(n130) );
  DFF_X1 reg_mem_reg_16__5_ ( .D(n6973), .CK(clk), .Q(n[2478]), .QN(n131) );
  DFF_X1 reg_mem_reg_16__4_ ( .D(n6972), .CK(clk), .Q(n[2477]), .QN(n132) );
  DFF_X1 reg_mem_reg_16__3_ ( .D(n6971), .CK(clk), .Q(n[2476]), .QN(n133) );
  DFF_X1 reg_mem_reg_16__2_ ( .D(n6970), .CK(clk), .Q(n[2475]), .QN(n134) );
  DFF_X1 reg_mem_reg_16__1_ ( .D(n6969), .CK(clk), .Q(n[2474]), .QN(n135) );
  DFF_X1 reg_mem_reg_16__0_ ( .D(n6968), .CK(clk), .Q(n[2473]), .QN(n136) );
  DFF_X1 reg_mem_reg_17__7_ ( .D(n6967), .CK(clk), .Q(n[2472]), .QN(n137) );
  DFF_X1 reg_mem_reg_17__6_ ( .D(n6966), .CK(clk), .Q(n[2471]), .QN(n138) );
  DFF_X1 reg_mem_reg_17__5_ ( .D(n6965), .CK(clk), .Q(n[2470]), .QN(n139) );
  DFF_X1 reg_mem_reg_17__4_ ( .D(n6964), .CK(clk), .Q(n[2469]), .QN(n140) );
  DFF_X1 reg_mem_reg_17__3_ ( .D(n6963), .CK(clk), .Q(n[2468]), .QN(n141) );
  DFF_X1 reg_mem_reg_17__2_ ( .D(n6962), .CK(clk), .Q(n[2467]), .QN(n142) );
  DFF_X1 reg_mem_reg_17__1_ ( .D(n6961), .CK(clk), .Q(n[2466]), .QN(n143) );
  DFF_X1 reg_mem_reg_17__0_ ( .D(n6960), .CK(clk), .Q(n[2465]), .QN(n144) );
  DFF_X1 reg_mem_reg_18__7_ ( .D(n6959), .CK(clk), .QN(n145) );
  DFF_X1 reg_mem_reg_18__6_ ( .D(n6958), .CK(clk), .QN(n146) );
  DFF_X1 reg_mem_reg_18__5_ ( .D(n6957), .CK(clk), .QN(n147) );
  DFF_X1 reg_mem_reg_18__4_ ( .D(n6956), .CK(clk), .QN(n148) );
  DFF_X1 reg_mem_reg_18__3_ ( .D(n6955), .CK(clk), .QN(n149) );
  DFF_X1 reg_mem_reg_18__2_ ( .D(n6954), .CK(clk), .QN(n150) );
  DFF_X1 reg_mem_reg_18__1_ ( .D(n6953), .CK(clk), .QN(n151) );
  DFF_X1 reg_mem_reg_18__0_ ( .D(n6952), .CK(clk), .QN(n152) );
  DFF_X1 reg_mem_reg_19__7_ ( .D(n6951), .CK(clk), .QN(n153) );
  DFF_X1 reg_mem_reg_19__6_ ( .D(n6950), .CK(clk), .QN(n154) );
  DFF_X1 reg_mem_reg_19__5_ ( .D(n6949), .CK(clk), .QN(n155) );
  DFF_X1 reg_mem_reg_19__4_ ( .D(n6948), .CK(clk), .QN(n156) );
  DFF_X1 reg_mem_reg_19__3_ ( .D(n6947), .CK(clk), .QN(n157) );
  DFF_X1 reg_mem_reg_19__2_ ( .D(n6946), .CK(clk), .QN(n158) );
  DFF_X1 reg_mem_reg_19__1_ ( .D(n6945), .CK(clk), .QN(n159) );
  DFF_X1 reg_mem_reg_19__0_ ( .D(n6944), .CK(clk), .QN(n160) );
  DFF_X1 reg_mem_reg_20__7_ ( .D(n6943), .CK(clk), .Q(n[2448]), .QN(n161) );
  DFF_X1 reg_mem_reg_20__6_ ( .D(n6942), .CK(clk), .Q(n[2447]), .QN(n162) );
  DFF_X1 reg_mem_reg_20__5_ ( .D(n6941), .CK(clk), .Q(n[2446]), .QN(n163) );
  DFF_X1 reg_mem_reg_20__4_ ( .D(n6940), .CK(clk), .Q(n[2445]), .QN(n164) );
  DFF_X1 reg_mem_reg_20__3_ ( .D(n6939), .CK(clk), .Q(n[2444]), .QN(n165) );
  DFF_X1 reg_mem_reg_20__2_ ( .D(n6938), .CK(clk), .Q(n[2443]), .QN(n166) );
  DFF_X1 reg_mem_reg_20__1_ ( .D(n6937), .CK(clk), .Q(n[2442]), .QN(n167) );
  DFF_X1 reg_mem_reg_20__0_ ( .D(n6936), .CK(clk), .Q(n[2441]), .QN(n168) );
  DFF_X1 reg_mem_reg_21__7_ ( .D(n6935), .CK(clk), .Q(n[2440]), .QN(n169) );
  DFF_X1 reg_mem_reg_21__6_ ( .D(n6934), .CK(clk), .Q(n[2439]), .QN(n170) );
  DFF_X1 reg_mem_reg_21__5_ ( .D(n6933), .CK(clk), .Q(n[2438]), .QN(n171) );
  DFF_X1 reg_mem_reg_21__4_ ( .D(n6932), .CK(clk), .Q(n[2437]), .QN(n172) );
  DFF_X1 reg_mem_reg_21__3_ ( .D(n6931), .CK(clk), .Q(n[2436]), .QN(n173) );
  DFF_X1 reg_mem_reg_21__2_ ( .D(n6930), .CK(clk), .Q(n[2435]), .QN(n174) );
  DFF_X1 reg_mem_reg_21__1_ ( .D(n6929), .CK(clk), .Q(n[2434]), .QN(n175) );
  DFF_X1 reg_mem_reg_21__0_ ( .D(n6928), .CK(clk), .Q(n[2433]), .QN(n176) );
  DFF_X1 reg_mem_reg_22__7_ ( .D(n6927), .CK(clk), .QN(n177) );
  DFF_X1 reg_mem_reg_22__6_ ( .D(n6926), .CK(clk), .QN(n178) );
  DFF_X1 reg_mem_reg_22__5_ ( .D(n6925), .CK(clk), .QN(n179) );
  DFF_X1 reg_mem_reg_22__4_ ( .D(n6924), .CK(clk), .QN(n180) );
  DFF_X1 reg_mem_reg_22__3_ ( .D(n6923), .CK(clk), .QN(n181) );
  DFF_X1 reg_mem_reg_22__2_ ( .D(n6922), .CK(clk), .QN(n182) );
  DFF_X1 reg_mem_reg_22__1_ ( .D(n6921), .CK(clk), .QN(n183) );
  DFF_X1 reg_mem_reg_22__0_ ( .D(n6920), .CK(clk), .QN(n184) );
  DFF_X1 reg_mem_reg_23__7_ ( .D(n6919), .CK(clk), .QN(n185) );
  DFF_X1 reg_mem_reg_23__6_ ( .D(n6918), .CK(clk), .QN(n186) );
  DFF_X1 reg_mem_reg_23__5_ ( .D(n6917), .CK(clk), .QN(n187) );
  DFF_X1 reg_mem_reg_23__4_ ( .D(n6916), .CK(clk), .QN(n188) );
  DFF_X1 reg_mem_reg_23__3_ ( .D(n6915), .CK(clk), .QN(n189) );
  DFF_X1 reg_mem_reg_23__2_ ( .D(n6914), .CK(clk), .QN(n190) );
  DFF_X1 reg_mem_reg_23__1_ ( .D(n6913), .CK(clk), .QN(n191) );
  DFF_X1 reg_mem_reg_23__0_ ( .D(n6912), .CK(clk), .QN(n192) );
  DFF_X1 reg_mem_reg_24__7_ ( .D(n6911), .CK(clk), .Q(n[2416]), .QN(n193) );
  DFF_X1 reg_mem_reg_24__6_ ( .D(n6910), .CK(clk), .Q(n[2415]), .QN(n194) );
  DFF_X1 reg_mem_reg_24__5_ ( .D(n6909), .CK(clk), .Q(n[2414]), .QN(n195) );
  DFF_X1 reg_mem_reg_24__4_ ( .D(n6908), .CK(clk), .Q(n[2413]), .QN(n196) );
  DFF_X1 reg_mem_reg_24__3_ ( .D(n6907), .CK(clk), .Q(n[2412]), .QN(n197) );
  DFF_X1 reg_mem_reg_24__2_ ( .D(n6906), .CK(clk), .Q(n[2411]), .QN(n198) );
  DFF_X1 reg_mem_reg_24__1_ ( .D(n6905), .CK(clk), .Q(n[2410]), .QN(n199) );
  DFF_X1 reg_mem_reg_24__0_ ( .D(n6904), .CK(clk), .Q(n[2409]), .QN(n200) );
  DFF_X1 reg_mem_reg_25__7_ ( .D(n6903), .CK(clk), .Q(n[2408]), .QN(n201) );
  DFF_X1 reg_mem_reg_25__6_ ( .D(n6902), .CK(clk), .Q(n[2407]), .QN(n202) );
  DFF_X1 reg_mem_reg_25__5_ ( .D(n6901), .CK(clk), .Q(n[2406]), .QN(n203) );
  DFF_X1 reg_mem_reg_25__4_ ( .D(n6900), .CK(clk), .Q(n[2405]), .QN(n204) );
  DFF_X1 reg_mem_reg_25__3_ ( .D(n6899), .CK(clk), .Q(n[2404]), .QN(n205) );
  DFF_X1 reg_mem_reg_25__2_ ( .D(n6898), .CK(clk), .Q(n[2403]), .QN(n206) );
  DFF_X1 reg_mem_reg_25__1_ ( .D(n6897), .CK(clk), .Q(n[2402]), .QN(n207) );
  DFF_X1 reg_mem_reg_25__0_ ( .D(n6896), .CK(clk), .Q(n[2401]), .QN(n208) );
  DFF_X1 reg_mem_reg_26__7_ ( .D(n6895), .CK(clk), .QN(n209) );
  DFF_X1 reg_mem_reg_26__6_ ( .D(n6894), .CK(clk), .QN(n210) );
  DFF_X1 reg_mem_reg_26__5_ ( .D(n6893), .CK(clk), .QN(n211) );
  DFF_X1 reg_mem_reg_26__4_ ( .D(n6892), .CK(clk), .QN(n212) );
  DFF_X1 reg_mem_reg_26__3_ ( .D(n6891), .CK(clk), .QN(n213) );
  DFF_X1 reg_mem_reg_26__2_ ( .D(n6890), .CK(clk), .QN(n214) );
  DFF_X1 reg_mem_reg_26__1_ ( .D(n6889), .CK(clk), .QN(n215) );
  DFF_X1 reg_mem_reg_26__0_ ( .D(n6888), .CK(clk), .QN(n216) );
  DFF_X1 reg_mem_reg_27__7_ ( .D(n6887), .CK(clk), .QN(n217) );
  DFF_X1 reg_mem_reg_27__6_ ( .D(n6886), .CK(clk), .QN(n218) );
  DFF_X1 reg_mem_reg_27__5_ ( .D(n6885), .CK(clk), .QN(n219) );
  DFF_X1 reg_mem_reg_27__4_ ( .D(n6884), .CK(clk), .QN(n220) );
  DFF_X1 reg_mem_reg_27__3_ ( .D(n6883), .CK(clk), .QN(n221) );
  DFF_X1 reg_mem_reg_27__2_ ( .D(n6882), .CK(clk), .QN(n222) );
  DFF_X1 reg_mem_reg_27__1_ ( .D(n6881), .CK(clk), .QN(n223) );
  DFF_X1 reg_mem_reg_27__0_ ( .D(n6880), .CK(clk), .QN(n224) );
  DFF_X1 reg_mem_reg_28__7_ ( .D(n6879), .CK(clk), .Q(n[2384]), .QN(n225) );
  DFF_X1 reg_mem_reg_28__6_ ( .D(n6878), .CK(clk), .Q(n[2383]), .QN(n226) );
  DFF_X1 reg_mem_reg_28__5_ ( .D(n6877), .CK(clk), .Q(n[2382]), .QN(n227) );
  DFF_X1 reg_mem_reg_28__4_ ( .D(n6876), .CK(clk), .Q(n[2381]), .QN(n228) );
  DFF_X1 reg_mem_reg_28__3_ ( .D(n6875), .CK(clk), .Q(n[2380]), .QN(n229) );
  DFF_X1 reg_mem_reg_28__2_ ( .D(n6874), .CK(clk), .Q(n[2379]), .QN(n230) );
  DFF_X1 reg_mem_reg_28__1_ ( .D(n6873), .CK(clk), .Q(n[2378]), .QN(n231) );
  DFF_X1 reg_mem_reg_28__0_ ( .D(n6872), .CK(clk), .Q(n[2377]), .QN(n232) );
  DFF_X1 reg_mem_reg_29__7_ ( .D(n6871), .CK(clk), .Q(n[2376]), .QN(n233) );
  DFF_X1 reg_mem_reg_29__6_ ( .D(n6870), .CK(clk), .Q(n[2375]), .QN(n234) );
  DFF_X1 reg_mem_reg_29__5_ ( .D(n6869), .CK(clk), .Q(n[2374]), .QN(n235) );
  DFF_X1 reg_mem_reg_29__4_ ( .D(n6868), .CK(clk), .Q(n[2373]), .QN(n236) );
  DFF_X1 reg_mem_reg_29__3_ ( .D(n6867), .CK(clk), .Q(n[2372]), .QN(n237) );
  DFF_X1 reg_mem_reg_29__2_ ( .D(n6866), .CK(clk), .Q(n[2371]), .QN(n238) );
  DFF_X1 reg_mem_reg_29__1_ ( .D(n6865), .CK(clk), .Q(n[2370]), .QN(n239) );
  DFF_X1 reg_mem_reg_29__0_ ( .D(n6864), .CK(clk), .Q(n[2369]), .QN(n240) );
  DFF_X1 reg_mem_reg_30__7_ ( .D(n6863), .CK(clk), .QN(n241) );
  DFF_X1 reg_mem_reg_30__6_ ( .D(n6862), .CK(clk), .QN(n242) );
  DFF_X1 reg_mem_reg_30__5_ ( .D(n6861), .CK(clk), .QN(n243) );
  DFF_X1 reg_mem_reg_30__4_ ( .D(n6860), .CK(clk), .QN(n244) );
  DFF_X1 reg_mem_reg_30__3_ ( .D(n6859), .CK(clk), .QN(n245) );
  DFF_X1 reg_mem_reg_30__2_ ( .D(n6858), .CK(clk), .QN(n246) );
  DFF_X1 reg_mem_reg_30__1_ ( .D(n6857), .CK(clk), .QN(n247) );
  DFF_X1 reg_mem_reg_30__0_ ( .D(n6856), .CK(clk), .QN(n248) );
  DFF_X1 reg_mem_reg_31__7_ ( .D(n6855), .CK(clk), .QN(n249) );
  DFF_X1 reg_mem_reg_31__6_ ( .D(n6854), .CK(clk), .QN(n250) );
  DFF_X1 reg_mem_reg_31__5_ ( .D(n6853), .CK(clk), .QN(n251) );
  DFF_X1 reg_mem_reg_31__4_ ( .D(n6852), .CK(clk), .QN(n252) );
  DFF_X1 reg_mem_reg_31__3_ ( .D(n6851), .CK(clk), .QN(n253) );
  DFF_X1 reg_mem_reg_31__2_ ( .D(n6850), .CK(clk), .QN(n254) );
  DFF_X1 reg_mem_reg_31__1_ ( .D(n6849), .CK(clk), .QN(n255) );
  DFF_X1 reg_mem_reg_31__0_ ( .D(n6848), .CK(clk), .QN(n256) );
  DFF_X1 reg_mem_reg_32__7_ ( .D(n6847), .CK(clk), .Q(n[2352]), .QN(n257) );
  DFF_X1 reg_mem_reg_32__6_ ( .D(n6846), .CK(clk), .Q(n[2351]), .QN(n258) );
  DFF_X1 reg_mem_reg_32__5_ ( .D(n6845), .CK(clk), .Q(n[2350]), .QN(n259) );
  DFF_X1 reg_mem_reg_32__4_ ( .D(n6844), .CK(clk), .Q(n[2349]), .QN(n260) );
  DFF_X1 reg_mem_reg_32__3_ ( .D(n6843), .CK(clk), .Q(n[2348]), .QN(n261) );
  DFF_X1 reg_mem_reg_32__2_ ( .D(n6842), .CK(clk), .Q(n[2347]), .QN(n262) );
  DFF_X1 reg_mem_reg_32__1_ ( .D(n6841), .CK(clk), .Q(n[2346]), .QN(n263) );
  DFF_X1 reg_mem_reg_32__0_ ( .D(n6840), .CK(clk), .Q(n[2345]), .QN(n264) );
  DFF_X1 reg_mem_reg_33__7_ ( .D(n6839), .CK(clk), .Q(n[2344]), .QN(n265) );
  DFF_X1 reg_mem_reg_33__6_ ( .D(n6838), .CK(clk), .Q(n[2343]), .QN(n266) );
  DFF_X1 reg_mem_reg_33__5_ ( .D(n6837), .CK(clk), .Q(n[2342]), .QN(n267) );
  DFF_X1 reg_mem_reg_33__4_ ( .D(n6836), .CK(clk), .Q(n[2341]), .QN(n268) );
  DFF_X1 reg_mem_reg_33__3_ ( .D(n6835), .CK(clk), .Q(n[2340]), .QN(n269) );
  DFF_X1 reg_mem_reg_33__2_ ( .D(n6834), .CK(clk), .Q(n[2339]), .QN(n270) );
  DFF_X1 reg_mem_reg_33__1_ ( .D(n6833), .CK(clk), .Q(n[2338]), .QN(n271) );
  DFF_X1 reg_mem_reg_33__0_ ( .D(n6832), .CK(clk), .Q(n[2337]), .QN(n272) );
  DFF_X1 reg_mem_reg_34__7_ ( .D(n6831), .CK(clk), .QN(n273) );
  DFF_X1 reg_mem_reg_34__6_ ( .D(n6830), .CK(clk), .QN(n274) );
  DFF_X1 reg_mem_reg_34__5_ ( .D(n6829), .CK(clk), .QN(n275) );
  DFF_X1 reg_mem_reg_34__4_ ( .D(n6828), .CK(clk), .QN(n276) );
  DFF_X1 reg_mem_reg_34__3_ ( .D(n6827), .CK(clk), .QN(n277) );
  DFF_X1 reg_mem_reg_34__2_ ( .D(n6826), .CK(clk), .QN(n278) );
  DFF_X1 reg_mem_reg_34__1_ ( .D(n6825), .CK(clk), .QN(n279) );
  DFF_X1 reg_mem_reg_34__0_ ( .D(n6824), .CK(clk), .QN(n280) );
  DFF_X1 reg_mem_reg_35__7_ ( .D(n6823), .CK(clk), .QN(n281) );
  DFF_X1 reg_mem_reg_35__6_ ( .D(n6822), .CK(clk), .QN(n282) );
  DFF_X1 reg_mem_reg_35__5_ ( .D(n6821), .CK(clk), .QN(n283) );
  DFF_X1 reg_mem_reg_35__4_ ( .D(n6820), .CK(clk), .QN(n284) );
  DFF_X1 reg_mem_reg_35__3_ ( .D(n6819), .CK(clk), .QN(n285) );
  DFF_X1 reg_mem_reg_35__2_ ( .D(n6818), .CK(clk), .QN(n286) );
  DFF_X1 reg_mem_reg_35__1_ ( .D(n6817), .CK(clk), .QN(n287) );
  DFF_X1 reg_mem_reg_35__0_ ( .D(n6816), .CK(clk), .QN(n288) );
  DFF_X1 reg_mem_reg_36__7_ ( .D(n6815), .CK(clk), .Q(n[2320]), .QN(n289) );
  DFF_X1 reg_mem_reg_36__6_ ( .D(n6814), .CK(clk), .Q(n[2319]), .QN(n290) );
  DFF_X1 reg_mem_reg_36__5_ ( .D(n6813), .CK(clk), .Q(n[2318]), .QN(n291) );
  DFF_X1 reg_mem_reg_36__4_ ( .D(n6812), .CK(clk), .Q(n[2317]), .QN(n292) );
  DFF_X1 reg_mem_reg_36__3_ ( .D(n6811), .CK(clk), .Q(n[2316]), .QN(n293) );
  DFF_X1 reg_mem_reg_36__2_ ( .D(n6810), .CK(clk), .Q(n[2315]), .QN(n294) );
  DFF_X1 reg_mem_reg_36__1_ ( .D(n6809), .CK(clk), .Q(n[2314]), .QN(n295) );
  DFF_X1 reg_mem_reg_36__0_ ( .D(n6808), .CK(clk), .Q(n[2313]), .QN(n296) );
  DFF_X1 reg_mem_reg_37__7_ ( .D(n6807), .CK(clk), .Q(n[2312]), .QN(n297) );
  DFF_X1 reg_mem_reg_37__6_ ( .D(n6806), .CK(clk), .Q(n[2311]), .QN(n298) );
  DFF_X1 reg_mem_reg_37__5_ ( .D(n6805), .CK(clk), .Q(n[2310]), .QN(n299) );
  DFF_X1 reg_mem_reg_37__4_ ( .D(n6804), .CK(clk), .Q(n[2309]), .QN(n300) );
  DFF_X1 reg_mem_reg_37__3_ ( .D(n6803), .CK(clk), .Q(n[2308]), .QN(n301) );
  DFF_X1 reg_mem_reg_37__2_ ( .D(n6802), .CK(clk), .Q(n[2307]), .QN(n302) );
  DFF_X1 reg_mem_reg_37__1_ ( .D(n6801), .CK(clk), .Q(n[2306]), .QN(n303) );
  DFF_X1 reg_mem_reg_37__0_ ( .D(n6800), .CK(clk), .Q(n[2305]), .QN(n304) );
  DFF_X1 reg_mem_reg_38__7_ ( .D(n6799), .CK(clk), .QN(n305) );
  DFF_X1 reg_mem_reg_38__6_ ( .D(n6798), .CK(clk), .QN(n306) );
  DFF_X1 reg_mem_reg_38__5_ ( .D(n6797), .CK(clk), .QN(n307) );
  DFF_X1 reg_mem_reg_38__4_ ( .D(n6796), .CK(clk), .QN(n308) );
  DFF_X1 reg_mem_reg_38__3_ ( .D(n6795), .CK(clk), .QN(n309) );
  DFF_X1 reg_mem_reg_38__2_ ( .D(n6794), .CK(clk), .QN(n310) );
  DFF_X1 reg_mem_reg_38__1_ ( .D(n6793), .CK(clk), .QN(n311) );
  DFF_X1 reg_mem_reg_38__0_ ( .D(n6792), .CK(clk), .QN(n312) );
  DFF_X1 reg_mem_reg_39__7_ ( .D(n6791), .CK(clk), .QN(n313) );
  DFF_X1 reg_mem_reg_39__6_ ( .D(n6790), .CK(clk), .QN(n314) );
  DFF_X1 reg_mem_reg_39__5_ ( .D(n6789), .CK(clk), .QN(n315) );
  DFF_X1 reg_mem_reg_39__4_ ( .D(n6788), .CK(clk), .QN(n316) );
  DFF_X1 reg_mem_reg_39__3_ ( .D(n6787), .CK(clk), .QN(n317) );
  DFF_X1 reg_mem_reg_39__2_ ( .D(n6786), .CK(clk), .QN(n318) );
  DFF_X1 reg_mem_reg_39__1_ ( .D(n6785), .CK(clk), .QN(n319) );
  DFF_X1 reg_mem_reg_39__0_ ( .D(n6784), .CK(clk), .QN(n320) );
  DFF_X1 reg_mem_reg_40__7_ ( .D(n6783), .CK(clk), .Q(n[2288]), .QN(n321) );
  DFF_X1 reg_mem_reg_40__6_ ( .D(n6782), .CK(clk), .Q(n[2287]), .QN(n322) );
  DFF_X1 reg_mem_reg_40__5_ ( .D(n6781), .CK(clk), .Q(n[2286]), .QN(n323) );
  DFF_X1 reg_mem_reg_40__4_ ( .D(n6780), .CK(clk), .Q(n[2285]), .QN(n324) );
  DFF_X1 reg_mem_reg_40__3_ ( .D(n6779), .CK(clk), .Q(n[2284]), .QN(n325) );
  DFF_X1 reg_mem_reg_40__2_ ( .D(n6778), .CK(clk), .Q(n[2283]), .QN(n326) );
  DFF_X1 reg_mem_reg_40__1_ ( .D(n6777), .CK(clk), .Q(n[2282]), .QN(n327) );
  DFF_X1 reg_mem_reg_40__0_ ( .D(n6776), .CK(clk), .Q(n[2281]), .QN(n328) );
  DFF_X1 reg_mem_reg_41__7_ ( .D(n6775), .CK(clk), .Q(n[2280]), .QN(n329) );
  DFF_X1 reg_mem_reg_41__6_ ( .D(n6774), .CK(clk), .Q(n[2279]), .QN(n330) );
  DFF_X1 reg_mem_reg_41__5_ ( .D(n6773), .CK(clk), .Q(n[2278]), .QN(n331) );
  DFF_X1 reg_mem_reg_41__4_ ( .D(n6772), .CK(clk), .Q(n[2277]), .QN(n332) );
  DFF_X1 reg_mem_reg_41__3_ ( .D(n6771), .CK(clk), .Q(n[2276]), .QN(n333) );
  DFF_X1 reg_mem_reg_41__2_ ( .D(n6770), .CK(clk), .Q(n[2275]), .QN(n334) );
  DFF_X1 reg_mem_reg_41__1_ ( .D(n6769), .CK(clk), .Q(n[2274]), .QN(n335) );
  DFF_X1 reg_mem_reg_41__0_ ( .D(n6768), .CK(clk), .Q(n[2273]), .QN(n336) );
  DFF_X1 reg_mem_reg_42__7_ ( .D(n6767), .CK(clk), .QN(n337) );
  DFF_X1 reg_mem_reg_42__6_ ( .D(n6766), .CK(clk), .QN(n338) );
  DFF_X1 reg_mem_reg_42__5_ ( .D(n6765), .CK(clk), .QN(n339) );
  DFF_X1 reg_mem_reg_42__4_ ( .D(n6764), .CK(clk), .QN(n340) );
  DFF_X1 reg_mem_reg_42__3_ ( .D(n6763), .CK(clk), .QN(n341) );
  DFF_X1 reg_mem_reg_42__2_ ( .D(n6762), .CK(clk), .QN(n342) );
  DFF_X1 reg_mem_reg_42__1_ ( .D(n6761), .CK(clk), .QN(n343) );
  DFF_X1 reg_mem_reg_42__0_ ( .D(n6760), .CK(clk), .QN(n344) );
  DFF_X1 reg_mem_reg_43__7_ ( .D(n6759), .CK(clk), .QN(n345) );
  DFF_X1 reg_mem_reg_43__6_ ( .D(n6758), .CK(clk), .QN(n346) );
  DFF_X1 reg_mem_reg_43__5_ ( .D(n6757), .CK(clk), .QN(n347) );
  DFF_X1 reg_mem_reg_43__4_ ( .D(n6756), .CK(clk), .QN(n348) );
  DFF_X1 reg_mem_reg_43__3_ ( .D(n6755), .CK(clk), .QN(n349) );
  DFF_X1 reg_mem_reg_43__2_ ( .D(n6754), .CK(clk), .QN(n350) );
  DFF_X1 reg_mem_reg_43__1_ ( .D(n6753), .CK(clk), .QN(n351) );
  DFF_X1 reg_mem_reg_43__0_ ( .D(n6752), .CK(clk), .QN(n352) );
  DFF_X1 reg_mem_reg_44__7_ ( .D(n6751), .CK(clk), .Q(n[2256]), .QN(n353) );
  DFF_X1 reg_mem_reg_44__6_ ( .D(n6750), .CK(clk), .Q(n[2255]), .QN(n354) );
  DFF_X1 reg_mem_reg_44__5_ ( .D(n6749), .CK(clk), .Q(n[2254]), .QN(n355) );
  DFF_X1 reg_mem_reg_44__4_ ( .D(n6748), .CK(clk), .Q(n[2253]), .QN(n356) );
  DFF_X1 reg_mem_reg_44__3_ ( .D(n6747), .CK(clk), .Q(n[2252]), .QN(n357) );
  DFF_X1 reg_mem_reg_44__2_ ( .D(n6746), .CK(clk), .Q(n[2251]), .QN(n358) );
  DFF_X1 reg_mem_reg_44__1_ ( .D(n6745), .CK(clk), .Q(n[2250]), .QN(n359) );
  DFF_X1 reg_mem_reg_44__0_ ( .D(n6744), .CK(clk), .Q(n[2249]), .QN(n360) );
  DFF_X1 reg_mem_reg_45__7_ ( .D(n6743), .CK(clk), .Q(n[2248]), .QN(n361) );
  DFF_X1 reg_mem_reg_45__6_ ( .D(n6742), .CK(clk), .Q(n[2247]), .QN(n362) );
  DFF_X1 reg_mem_reg_45__5_ ( .D(n6741), .CK(clk), .Q(n[2246]), .QN(n363) );
  DFF_X1 reg_mem_reg_45__4_ ( .D(n6740), .CK(clk), .Q(n[2245]), .QN(n364) );
  DFF_X1 reg_mem_reg_45__3_ ( .D(n6739), .CK(clk), .Q(n[2244]), .QN(n365) );
  DFF_X1 reg_mem_reg_45__2_ ( .D(n6738), .CK(clk), .Q(n[2243]), .QN(n366) );
  DFF_X1 reg_mem_reg_45__1_ ( .D(n6737), .CK(clk), .Q(n[2242]), .QN(n367) );
  DFF_X1 reg_mem_reg_45__0_ ( .D(n6736), .CK(clk), .Q(n[2241]), .QN(n368) );
  DFF_X1 reg_mem_reg_46__7_ ( .D(n6735), .CK(clk), .QN(n369) );
  DFF_X1 reg_mem_reg_46__6_ ( .D(n6734), .CK(clk), .QN(n370) );
  DFF_X1 reg_mem_reg_46__5_ ( .D(n6733), .CK(clk), .QN(n371) );
  DFF_X1 reg_mem_reg_46__4_ ( .D(n6732), .CK(clk), .QN(n372) );
  DFF_X1 reg_mem_reg_46__3_ ( .D(n6731), .CK(clk), .QN(n373) );
  DFF_X1 reg_mem_reg_46__2_ ( .D(n6730), .CK(clk), .QN(n374) );
  DFF_X1 reg_mem_reg_46__1_ ( .D(n6729), .CK(clk), .QN(n375) );
  DFF_X1 reg_mem_reg_46__0_ ( .D(n6728), .CK(clk), .QN(n376) );
  DFF_X1 reg_mem_reg_47__7_ ( .D(n6727), .CK(clk), .QN(n377) );
  DFF_X1 reg_mem_reg_47__6_ ( .D(n6726), .CK(clk), .QN(n378) );
  DFF_X1 reg_mem_reg_47__5_ ( .D(n6725), .CK(clk), .QN(n379) );
  DFF_X1 reg_mem_reg_47__4_ ( .D(n6724), .CK(clk), .QN(n380) );
  DFF_X1 reg_mem_reg_47__3_ ( .D(n6723), .CK(clk), .QN(n381) );
  DFF_X1 reg_mem_reg_47__2_ ( .D(n6722), .CK(clk), .QN(n382) );
  DFF_X1 reg_mem_reg_47__1_ ( .D(n6721), .CK(clk), .QN(n383) );
  DFF_X1 reg_mem_reg_47__0_ ( .D(n6720), .CK(clk), .QN(n384) );
  DFF_X1 reg_mem_reg_48__7_ ( .D(n6719), .CK(clk), .Q(n[2224]), .QN(n385) );
  DFF_X1 reg_mem_reg_48__6_ ( .D(n6718), .CK(clk), .Q(n[2223]), .QN(n386) );
  DFF_X1 reg_mem_reg_48__5_ ( .D(n6717), .CK(clk), .Q(n[2222]), .QN(n387) );
  DFF_X1 reg_mem_reg_48__4_ ( .D(n6716), .CK(clk), .Q(n[2221]), .QN(n388) );
  DFF_X1 reg_mem_reg_48__3_ ( .D(n6715), .CK(clk), .Q(n[2220]), .QN(n389) );
  DFF_X1 reg_mem_reg_48__2_ ( .D(n6714), .CK(clk), .Q(n[2219]), .QN(n390) );
  DFF_X1 reg_mem_reg_48__1_ ( .D(n6713), .CK(clk), .Q(n[2218]), .QN(n391) );
  DFF_X1 reg_mem_reg_48__0_ ( .D(n6712), .CK(clk), .Q(n[2217]), .QN(n392) );
  DFF_X1 reg_mem_reg_49__7_ ( .D(n6711), .CK(clk), .Q(n[2216]), .QN(n393) );
  DFF_X1 reg_mem_reg_49__6_ ( .D(n6710), .CK(clk), .Q(n[2215]), .QN(n394) );
  DFF_X1 reg_mem_reg_49__5_ ( .D(n6709), .CK(clk), .Q(n[2214]), .QN(n395) );
  DFF_X1 reg_mem_reg_49__4_ ( .D(n6708), .CK(clk), .Q(n[2213]), .QN(n396) );
  DFF_X1 reg_mem_reg_49__3_ ( .D(n6707), .CK(clk), .Q(n[2212]), .QN(n397) );
  DFF_X1 reg_mem_reg_49__2_ ( .D(n6706), .CK(clk), .Q(n[2211]), .QN(n398) );
  DFF_X1 reg_mem_reg_49__1_ ( .D(n6705), .CK(clk), .Q(n[2210]), .QN(n399) );
  DFF_X1 reg_mem_reg_49__0_ ( .D(n6704), .CK(clk), .Q(n[2209]), .QN(n400) );
  DFF_X1 reg_mem_reg_50__7_ ( .D(n6703), .CK(clk), .QN(n401) );
  DFF_X1 reg_mem_reg_50__6_ ( .D(n6702), .CK(clk), .QN(n402) );
  DFF_X1 reg_mem_reg_50__5_ ( .D(n6701), .CK(clk), .QN(n403) );
  DFF_X1 reg_mem_reg_50__4_ ( .D(n6700), .CK(clk), .QN(n404) );
  DFF_X1 reg_mem_reg_50__3_ ( .D(n6699), .CK(clk), .QN(n405) );
  DFF_X1 reg_mem_reg_50__2_ ( .D(n6698), .CK(clk), .QN(n406) );
  DFF_X1 reg_mem_reg_50__1_ ( .D(n6697), .CK(clk), .QN(n407) );
  DFF_X1 reg_mem_reg_50__0_ ( .D(n6696), .CK(clk), .QN(n408) );
  DFF_X1 reg_mem_reg_51__7_ ( .D(n6695), .CK(clk), .QN(n409) );
  DFF_X1 reg_mem_reg_51__6_ ( .D(n6694), .CK(clk), .QN(n410) );
  DFF_X1 reg_mem_reg_51__5_ ( .D(n6693), .CK(clk), .QN(n411) );
  DFF_X1 reg_mem_reg_51__4_ ( .D(n6692), .CK(clk), .QN(n412) );
  DFF_X1 reg_mem_reg_51__3_ ( .D(n6691), .CK(clk), .QN(n413) );
  DFF_X1 reg_mem_reg_51__2_ ( .D(n6690), .CK(clk), .QN(n414) );
  DFF_X1 reg_mem_reg_51__1_ ( .D(n6689), .CK(clk), .QN(n415) );
  DFF_X1 reg_mem_reg_51__0_ ( .D(n6688), .CK(clk), .QN(n416) );
  DFF_X1 reg_mem_reg_52__7_ ( .D(n6687), .CK(clk), .Q(n[2192]), .QN(n417) );
  DFF_X1 reg_mem_reg_52__6_ ( .D(n6686), .CK(clk), .Q(n[2191]), .QN(n418) );
  DFF_X1 reg_mem_reg_52__5_ ( .D(n6685), .CK(clk), .Q(n[2190]), .QN(n419) );
  DFF_X1 reg_mem_reg_52__4_ ( .D(n6684), .CK(clk), .Q(n[2189]), .QN(n420) );
  DFF_X1 reg_mem_reg_52__3_ ( .D(n6683), .CK(clk), .Q(n[2188]), .QN(n421) );
  DFF_X1 reg_mem_reg_52__2_ ( .D(n6682), .CK(clk), .Q(n[2187]), .QN(n422) );
  DFF_X1 reg_mem_reg_52__1_ ( .D(n6681), .CK(clk), .Q(n[2186]), .QN(n423) );
  DFF_X1 reg_mem_reg_52__0_ ( .D(n6680), .CK(clk), .Q(n[2185]), .QN(n424) );
  DFF_X1 reg_mem_reg_53__7_ ( .D(n6679), .CK(clk), .Q(n[2184]), .QN(n425) );
  DFF_X1 reg_mem_reg_53__6_ ( .D(n6678), .CK(clk), .Q(n[2183]), .QN(n426) );
  DFF_X1 reg_mem_reg_53__5_ ( .D(n6677), .CK(clk), .Q(n[2182]), .QN(n427) );
  DFF_X1 reg_mem_reg_53__4_ ( .D(n6676), .CK(clk), .Q(n[2181]), .QN(n428) );
  DFF_X1 reg_mem_reg_53__3_ ( .D(n6675), .CK(clk), .Q(n[2180]), .QN(n429) );
  DFF_X1 reg_mem_reg_53__2_ ( .D(n6674), .CK(clk), .Q(n[2179]), .QN(n430) );
  DFF_X1 reg_mem_reg_53__1_ ( .D(n6673), .CK(clk), .Q(n[2178]), .QN(n431) );
  DFF_X1 reg_mem_reg_53__0_ ( .D(n6672), .CK(clk), .Q(n[2177]), .QN(n432) );
  DFF_X1 reg_mem_reg_54__7_ ( .D(n6671), .CK(clk), .QN(n433) );
  DFF_X1 reg_mem_reg_54__6_ ( .D(n6670), .CK(clk), .QN(n434) );
  DFF_X1 reg_mem_reg_54__5_ ( .D(n6669), .CK(clk), .QN(n435) );
  DFF_X1 reg_mem_reg_54__4_ ( .D(n6668), .CK(clk), .QN(n436) );
  DFF_X1 reg_mem_reg_54__3_ ( .D(n6667), .CK(clk), .QN(n437) );
  DFF_X1 reg_mem_reg_54__2_ ( .D(n6666), .CK(clk), .QN(n438) );
  DFF_X1 reg_mem_reg_54__1_ ( .D(n6665), .CK(clk), .QN(n439) );
  DFF_X1 reg_mem_reg_54__0_ ( .D(n6664), .CK(clk), .QN(n440) );
  DFF_X1 reg_mem_reg_55__7_ ( .D(n6663), .CK(clk), .QN(n441) );
  DFF_X1 reg_mem_reg_55__6_ ( .D(n6662), .CK(clk), .QN(n442) );
  DFF_X1 reg_mem_reg_55__5_ ( .D(n6661), .CK(clk), .QN(n443) );
  DFF_X1 reg_mem_reg_55__4_ ( .D(n6660), .CK(clk), .QN(n444) );
  DFF_X1 reg_mem_reg_55__3_ ( .D(n6659), .CK(clk), .QN(n445) );
  DFF_X1 reg_mem_reg_55__2_ ( .D(n6658), .CK(clk), .QN(n446) );
  DFF_X1 reg_mem_reg_55__1_ ( .D(n6657), .CK(clk), .QN(n447) );
  DFF_X1 reg_mem_reg_55__0_ ( .D(n6656), .CK(clk), .QN(n448) );
  DFF_X1 reg_mem_reg_56__7_ ( .D(n6655), .CK(clk), .Q(n[2160]), .QN(n449) );
  DFF_X1 reg_mem_reg_56__6_ ( .D(n6654), .CK(clk), .Q(n[2159]), .QN(n450) );
  DFF_X1 reg_mem_reg_56__5_ ( .D(n6653), .CK(clk), .Q(n[2158]), .QN(n451) );
  DFF_X1 reg_mem_reg_56__4_ ( .D(n6652), .CK(clk), .Q(n[2157]), .QN(n452) );
  DFF_X1 reg_mem_reg_56__3_ ( .D(n6651), .CK(clk), .Q(n[2156]), .QN(n453) );
  DFF_X1 reg_mem_reg_56__2_ ( .D(n6650), .CK(clk), .Q(n[2155]), .QN(n454) );
  DFF_X1 reg_mem_reg_56__1_ ( .D(n6649), .CK(clk), .Q(n[2154]), .QN(n455) );
  DFF_X1 reg_mem_reg_56__0_ ( .D(n6648), .CK(clk), .Q(n[2153]), .QN(n456) );
  DFF_X1 reg_mem_reg_57__7_ ( .D(n6647), .CK(clk), .Q(n[2152]), .QN(n457) );
  DFF_X1 reg_mem_reg_57__6_ ( .D(n6646), .CK(clk), .Q(n[2151]), .QN(n458) );
  DFF_X1 reg_mem_reg_57__5_ ( .D(n6645), .CK(clk), .Q(n[2150]), .QN(n459) );
  DFF_X1 reg_mem_reg_57__4_ ( .D(n6644), .CK(clk), .Q(n[2149]), .QN(n460) );
  DFF_X1 reg_mem_reg_57__3_ ( .D(n6643), .CK(clk), .Q(n[2148]), .QN(n461) );
  DFF_X1 reg_mem_reg_57__2_ ( .D(n6642), .CK(clk), .Q(n[2147]), .QN(n462) );
  DFF_X1 reg_mem_reg_57__1_ ( .D(n6641), .CK(clk), .Q(n[2146]), .QN(n463) );
  DFF_X1 reg_mem_reg_57__0_ ( .D(n6640), .CK(clk), .Q(n[2145]), .QN(n464) );
  DFF_X1 reg_mem_reg_58__7_ ( .D(n6639), .CK(clk), .QN(n465) );
  DFF_X1 reg_mem_reg_58__6_ ( .D(n6638), .CK(clk), .QN(n466) );
  DFF_X1 reg_mem_reg_58__5_ ( .D(n6637), .CK(clk), .QN(n467) );
  DFF_X1 reg_mem_reg_58__4_ ( .D(n6636), .CK(clk), .QN(n468) );
  DFF_X1 reg_mem_reg_58__3_ ( .D(n6635), .CK(clk), .QN(n469) );
  DFF_X1 reg_mem_reg_58__2_ ( .D(n6634), .CK(clk), .QN(n470) );
  DFF_X1 reg_mem_reg_58__1_ ( .D(n6633), .CK(clk), .QN(n471) );
  DFF_X1 reg_mem_reg_58__0_ ( .D(n6632), .CK(clk), .QN(n472) );
  DFF_X1 reg_mem_reg_59__7_ ( .D(n6631), .CK(clk), .QN(n473) );
  DFF_X1 reg_mem_reg_59__6_ ( .D(n6630), .CK(clk), .QN(n474) );
  DFF_X1 reg_mem_reg_59__5_ ( .D(n6629), .CK(clk), .QN(n475) );
  DFF_X1 reg_mem_reg_59__4_ ( .D(n6628), .CK(clk), .QN(n476) );
  DFF_X1 reg_mem_reg_59__3_ ( .D(n6627), .CK(clk), .QN(n477) );
  DFF_X1 reg_mem_reg_59__2_ ( .D(n6626), .CK(clk), .QN(n478) );
  DFF_X1 reg_mem_reg_59__1_ ( .D(n6625), .CK(clk), .QN(n479) );
  DFF_X1 reg_mem_reg_59__0_ ( .D(n6624), .CK(clk), .QN(n480) );
  DFF_X1 reg_mem_reg_60__7_ ( .D(n6623), .CK(clk), .Q(n[2128]), .QN(n481) );
  DFF_X1 reg_mem_reg_60__6_ ( .D(n6622), .CK(clk), .Q(n[2127]), .QN(n482) );
  DFF_X1 reg_mem_reg_60__5_ ( .D(n6621), .CK(clk), .Q(n[2126]), .QN(n483) );
  DFF_X1 reg_mem_reg_60__4_ ( .D(n6620), .CK(clk), .Q(n[2125]), .QN(n484) );
  DFF_X1 reg_mem_reg_60__3_ ( .D(n6619), .CK(clk), .Q(n[2124]), .QN(n485) );
  DFF_X1 reg_mem_reg_60__2_ ( .D(n6618), .CK(clk), .Q(n[2123]), .QN(n486) );
  DFF_X1 reg_mem_reg_60__1_ ( .D(n6617), .CK(clk), .Q(n[2122]), .QN(n487) );
  DFF_X1 reg_mem_reg_60__0_ ( .D(n6616), .CK(clk), .Q(n[2121]), .QN(n488) );
  DFF_X1 reg_mem_reg_61__7_ ( .D(n6615), .CK(clk), .Q(n[2120]), .QN(n489) );
  DFF_X1 reg_mem_reg_61__6_ ( .D(n6614), .CK(clk), .Q(n[2119]), .QN(n490) );
  DFF_X1 reg_mem_reg_61__5_ ( .D(n6613), .CK(clk), .Q(n[2118]), .QN(n491) );
  DFF_X1 reg_mem_reg_61__4_ ( .D(n6612), .CK(clk), .Q(n[2117]), .QN(n492) );
  DFF_X1 reg_mem_reg_61__3_ ( .D(n6611), .CK(clk), .Q(n[2116]), .QN(n493) );
  DFF_X1 reg_mem_reg_61__2_ ( .D(n6610), .CK(clk), .Q(n[2115]), .QN(n494) );
  DFF_X1 reg_mem_reg_61__1_ ( .D(n6609), .CK(clk), .Q(n[2114]), .QN(n495) );
  DFF_X1 reg_mem_reg_61__0_ ( .D(n6608), .CK(clk), .Q(n[2113]), .QN(n496) );
  DFF_X1 reg_mem_reg_62__7_ ( .D(n6607), .CK(clk), .QN(n497) );
  DFF_X1 reg_mem_reg_62__6_ ( .D(n6606), .CK(clk), .QN(n498) );
  DFF_X1 reg_mem_reg_62__5_ ( .D(n6605), .CK(clk), .QN(n499) );
  DFF_X1 reg_mem_reg_62__4_ ( .D(n6604), .CK(clk), .QN(n500) );
  DFF_X1 reg_mem_reg_62__3_ ( .D(n6603), .CK(clk), .QN(n501) );
  DFF_X1 reg_mem_reg_62__2_ ( .D(n6602), .CK(clk), .QN(n502) );
  DFF_X1 reg_mem_reg_62__1_ ( .D(n6601), .CK(clk), .QN(n503) );
  DFF_X1 reg_mem_reg_62__0_ ( .D(n6600), .CK(clk), .QN(n504) );
  DFF_X1 reg_mem_reg_63__7_ ( .D(n6599), .CK(clk), .QN(n505) );
  DFF_X1 reg_mem_reg_63__6_ ( .D(n6598), .CK(clk), .QN(n506) );
  DFF_X1 reg_mem_reg_63__5_ ( .D(n6597), .CK(clk), .QN(n507) );
  DFF_X1 reg_mem_reg_63__4_ ( .D(n6596), .CK(clk), .QN(n508) );
  DFF_X1 reg_mem_reg_63__3_ ( .D(n6595), .CK(clk), .QN(n509) );
  DFF_X1 reg_mem_reg_63__2_ ( .D(n6594), .CK(clk), .QN(n510) );
  DFF_X1 reg_mem_reg_63__1_ ( .D(n6593), .CK(clk), .QN(n511) );
  DFF_X1 reg_mem_reg_63__0_ ( .D(n6592), .CK(clk), .QN(n512) );
  DFF_X1 reg_mem_reg_64__7_ ( .D(n6591), .CK(clk), .Q(n[2096]), .QN(n513) );
  DFF_X1 reg_mem_reg_64__6_ ( .D(n6590), .CK(clk), .Q(n[2095]), .QN(n514) );
  DFF_X1 reg_mem_reg_64__5_ ( .D(n6589), .CK(clk), .Q(n[2094]), .QN(n515) );
  DFF_X1 reg_mem_reg_64__4_ ( .D(n6588), .CK(clk), .Q(n[2093]), .QN(n516) );
  DFF_X1 reg_mem_reg_64__3_ ( .D(n6587), .CK(clk), .Q(n[2092]), .QN(n517) );
  DFF_X1 reg_mem_reg_64__2_ ( .D(n6586), .CK(clk), .Q(n[2091]), .QN(n518) );
  DFF_X1 reg_mem_reg_64__1_ ( .D(n6585), .CK(clk), .Q(n[2090]), .QN(n519) );
  DFF_X1 reg_mem_reg_64__0_ ( .D(n6584), .CK(clk), .Q(n[2089]), .QN(n520) );
  DFF_X1 reg_mem_reg_65__7_ ( .D(n6583), .CK(clk), .Q(n[2088]), .QN(n521) );
  DFF_X1 reg_mem_reg_65__6_ ( .D(n6582), .CK(clk), .Q(n[2087]), .QN(n522) );
  DFF_X1 reg_mem_reg_65__5_ ( .D(n6581), .CK(clk), .Q(n[2086]), .QN(n523) );
  DFF_X1 reg_mem_reg_65__4_ ( .D(n6580), .CK(clk), .Q(n[2085]), .QN(n524) );
  DFF_X1 reg_mem_reg_65__3_ ( .D(n6579), .CK(clk), .Q(n[2084]), .QN(n525) );
  DFF_X1 reg_mem_reg_65__2_ ( .D(n6578), .CK(clk), .Q(n[2083]), .QN(n526) );
  DFF_X1 reg_mem_reg_65__1_ ( .D(n6577), .CK(clk), .Q(n[2082]), .QN(n527) );
  DFF_X1 reg_mem_reg_65__0_ ( .D(n6576), .CK(clk), .Q(n[2081]), .QN(n528) );
  DFF_X1 reg_mem_reg_66__7_ ( .D(n6575), .CK(clk), .QN(n529) );
  DFF_X1 reg_mem_reg_66__6_ ( .D(n6574), .CK(clk), .QN(n530) );
  DFF_X1 reg_mem_reg_66__5_ ( .D(n6573), .CK(clk), .QN(n531) );
  DFF_X1 reg_mem_reg_66__4_ ( .D(n6572), .CK(clk), .QN(n532) );
  DFF_X1 reg_mem_reg_66__3_ ( .D(n6571), .CK(clk), .QN(n533) );
  DFF_X1 reg_mem_reg_66__2_ ( .D(n6570), .CK(clk), .QN(n534) );
  DFF_X1 reg_mem_reg_66__1_ ( .D(n6569), .CK(clk), .QN(n535) );
  DFF_X1 reg_mem_reg_66__0_ ( .D(n6568), .CK(clk), .QN(n536) );
  DFF_X1 reg_mem_reg_67__7_ ( .D(n6567), .CK(clk), .QN(n537) );
  DFF_X1 reg_mem_reg_67__6_ ( .D(n6566), .CK(clk), .QN(n538) );
  DFF_X1 reg_mem_reg_67__5_ ( .D(n6565), .CK(clk), .QN(n539) );
  DFF_X1 reg_mem_reg_67__4_ ( .D(n6564), .CK(clk), .QN(n540) );
  DFF_X1 reg_mem_reg_67__3_ ( .D(n6563), .CK(clk), .QN(n541) );
  DFF_X1 reg_mem_reg_67__2_ ( .D(n6562), .CK(clk), .QN(n542) );
  DFF_X1 reg_mem_reg_67__1_ ( .D(n6561), .CK(clk), .QN(n543) );
  DFF_X1 reg_mem_reg_67__0_ ( .D(n6560), .CK(clk), .QN(n544) );
  DFF_X1 reg_mem_reg_68__7_ ( .D(n6559), .CK(clk), .Q(n[2064]), .QN(n545) );
  DFF_X1 reg_mem_reg_68__6_ ( .D(n6558), .CK(clk), .Q(n[2063]), .QN(n546) );
  DFF_X1 reg_mem_reg_68__5_ ( .D(n6557), .CK(clk), .Q(n[2062]), .QN(n547) );
  DFF_X1 reg_mem_reg_68__4_ ( .D(n6556), .CK(clk), .Q(n[2061]), .QN(n548) );
  DFF_X1 reg_mem_reg_68__3_ ( .D(n6555), .CK(clk), .Q(n[2060]), .QN(n549) );
  DFF_X1 reg_mem_reg_68__2_ ( .D(n6554), .CK(clk), .Q(n[2059]), .QN(n550) );
  DFF_X1 reg_mem_reg_68__1_ ( .D(n6553), .CK(clk), .Q(n[2058]), .QN(n551) );
  DFF_X1 reg_mem_reg_68__0_ ( .D(n6552), .CK(clk), .Q(n[2057]), .QN(n552) );
  DFF_X1 reg_mem_reg_69__7_ ( .D(n6551), .CK(clk), .Q(n[2056]), .QN(n553) );
  DFF_X1 reg_mem_reg_69__6_ ( .D(n6550), .CK(clk), .Q(n[2055]), .QN(n554) );
  DFF_X1 reg_mem_reg_69__5_ ( .D(n6549), .CK(clk), .Q(n[2054]), .QN(n555) );
  DFF_X1 reg_mem_reg_69__4_ ( .D(n6548), .CK(clk), .Q(n[2053]), .QN(n556) );
  DFF_X1 reg_mem_reg_69__3_ ( .D(n6547), .CK(clk), .Q(n[2052]), .QN(n557) );
  DFF_X1 reg_mem_reg_69__2_ ( .D(n6546), .CK(clk), .Q(n[2051]), .QN(n558) );
  DFF_X1 reg_mem_reg_69__1_ ( .D(n6545), .CK(clk), .Q(n[2050]), .QN(n559) );
  DFF_X1 reg_mem_reg_69__0_ ( .D(n6544), .CK(clk), .Q(n[2049]), .QN(n560) );
  DFF_X1 reg_mem_reg_70__7_ ( .D(n6543), .CK(clk), .QN(n561) );
  DFF_X1 reg_mem_reg_70__6_ ( .D(n6542), .CK(clk), .QN(n562) );
  DFF_X1 reg_mem_reg_70__5_ ( .D(n6541), .CK(clk), .QN(n563) );
  DFF_X1 reg_mem_reg_70__4_ ( .D(n6540), .CK(clk), .QN(n564) );
  DFF_X1 reg_mem_reg_70__3_ ( .D(n6539), .CK(clk), .QN(n565) );
  DFF_X1 reg_mem_reg_70__2_ ( .D(n6538), .CK(clk), .QN(n566) );
  DFF_X1 reg_mem_reg_70__1_ ( .D(n6537), .CK(clk), .QN(n567) );
  DFF_X1 reg_mem_reg_70__0_ ( .D(n6536), .CK(clk), .QN(n568) );
  DFF_X1 reg_mem_reg_71__7_ ( .D(n6535), .CK(clk), .QN(n569) );
  DFF_X1 reg_mem_reg_71__6_ ( .D(n6534), .CK(clk), .QN(n570) );
  DFF_X1 reg_mem_reg_71__5_ ( .D(n6533), .CK(clk), .QN(n571) );
  DFF_X1 reg_mem_reg_71__4_ ( .D(n6532), .CK(clk), .QN(n572) );
  DFF_X1 reg_mem_reg_71__3_ ( .D(n6531), .CK(clk), .QN(n573) );
  DFF_X1 reg_mem_reg_71__2_ ( .D(n6530), .CK(clk), .QN(n574) );
  DFF_X1 reg_mem_reg_71__1_ ( .D(n6529), .CK(clk), .QN(n575) );
  DFF_X1 reg_mem_reg_71__0_ ( .D(n6528), .CK(clk), .QN(n576) );
  DFF_X1 reg_mem_reg_72__7_ ( .D(n6527), .CK(clk), .Q(n[2032]), .QN(n593) );
  DFF_X1 reg_mem_reg_72__6_ ( .D(n6526), .CK(clk), .Q(n[2031]), .QN(n594) );
  DFF_X1 reg_mem_reg_72__5_ ( .D(n6525), .CK(clk), .Q(n[2030]), .QN(n595) );
  DFF_X1 reg_mem_reg_72__4_ ( .D(n6524), .CK(clk), .Q(n[2029]), .QN(n596) );
  DFF_X1 reg_mem_reg_72__3_ ( .D(n6523), .CK(clk), .Q(n[2028]), .QN(n597) );
  DFF_X1 reg_mem_reg_72__2_ ( .D(n6522), .CK(clk), .Q(n[2027]), .QN(n598) );
  DFF_X1 reg_mem_reg_72__1_ ( .D(n6521), .CK(clk), .Q(n[2026]), .QN(n599) );
  DFF_X1 reg_mem_reg_72__0_ ( .D(n6520), .CK(clk), .Q(n[2025]), .QN(n600) );
  DFF_X1 reg_mem_reg_73__7_ ( .D(n6519), .CK(clk), .Q(n[2024]), .QN(n601) );
  DFF_X1 reg_mem_reg_73__6_ ( .D(n6518), .CK(clk), .Q(n[2023]), .QN(n602) );
  DFF_X1 reg_mem_reg_73__5_ ( .D(n6517), .CK(clk), .Q(n[2022]), .QN(n603) );
  DFF_X1 reg_mem_reg_73__4_ ( .D(n6516), .CK(clk), .Q(n[2021]), .QN(n604) );
  DFF_X1 reg_mem_reg_73__3_ ( .D(n6515), .CK(clk), .Q(n[2020]), .QN(n605) );
  DFF_X1 reg_mem_reg_73__2_ ( .D(n6514), .CK(clk), .Q(n[2019]), .QN(n606) );
  DFF_X1 reg_mem_reg_73__1_ ( .D(n6513), .CK(clk), .Q(n[2018]), .QN(n607) );
  DFF_X1 reg_mem_reg_73__0_ ( .D(n6512), .CK(clk), .Q(n[2017]), .QN(n608) );
  DFF_X1 reg_mem_reg_74__7_ ( .D(n6511), .CK(clk), .QN(n625) );
  DFF_X1 reg_mem_reg_74__6_ ( .D(n6510), .CK(clk), .QN(n626) );
  DFF_X1 reg_mem_reg_74__5_ ( .D(n6509), .CK(clk), .QN(n627) );
  DFF_X1 reg_mem_reg_74__4_ ( .D(n6508), .CK(clk), .QN(n628) );
  DFF_X1 reg_mem_reg_74__3_ ( .D(n6507), .CK(clk), .QN(n629) );
  DFF_X1 reg_mem_reg_74__2_ ( .D(n6506), .CK(clk), .QN(n630) );
  DFF_X1 reg_mem_reg_74__1_ ( .D(n6505), .CK(clk), .QN(n631) );
  DFF_X1 reg_mem_reg_74__0_ ( .D(n6504), .CK(clk), .QN(n632) );
  DFF_X1 reg_mem_reg_75__7_ ( .D(n6503), .CK(clk), .QN(n633) );
  DFF_X1 reg_mem_reg_75__6_ ( .D(n6502), .CK(clk), .QN(n634) );
  DFF_X1 reg_mem_reg_75__5_ ( .D(n6501), .CK(clk), .QN(n635) );
  DFF_X1 reg_mem_reg_75__4_ ( .D(n6500), .CK(clk), .QN(n636) );
  DFF_X1 reg_mem_reg_75__3_ ( .D(n6499), .CK(clk), .QN(n637) );
  DFF_X1 reg_mem_reg_75__2_ ( .D(n6498), .CK(clk), .QN(n638) );
  DFF_X1 reg_mem_reg_75__1_ ( .D(n6497), .CK(clk), .QN(n639) );
  DFF_X1 reg_mem_reg_75__0_ ( .D(n6496), .CK(clk), .QN(n640) );
  DFF_X1 reg_mem_reg_76__7_ ( .D(n6495), .CK(clk), .Q(n[2000]), .QN(n657) );
  DFF_X1 reg_mem_reg_76__6_ ( .D(n6494), .CK(clk), .Q(n[1999]), .QN(n658) );
  DFF_X1 reg_mem_reg_76__5_ ( .D(n6493), .CK(clk), .Q(n[1998]), .QN(n659) );
  DFF_X1 reg_mem_reg_76__4_ ( .D(n6492), .CK(clk), .Q(n[1997]), .QN(n660) );
  DFF_X1 reg_mem_reg_76__3_ ( .D(n6491), .CK(clk), .Q(n[1996]), .QN(n661) );
  DFF_X1 reg_mem_reg_76__2_ ( .D(n6490), .CK(clk), .Q(n[1995]), .QN(n662) );
  DFF_X1 reg_mem_reg_76__1_ ( .D(n6489), .CK(clk), .Q(n[1994]), .QN(n663) );
  DFF_X1 reg_mem_reg_76__0_ ( .D(n6488), .CK(clk), .Q(n[1993]), .QN(n664) );
  DFF_X1 reg_mem_reg_77__7_ ( .D(n6487), .CK(clk), .Q(n[1992]), .QN(n665) );
  DFF_X1 reg_mem_reg_77__6_ ( .D(n6486), .CK(clk), .Q(n[1991]), .QN(n666) );
  DFF_X1 reg_mem_reg_77__5_ ( .D(n6485), .CK(clk), .Q(n[1990]), .QN(n667) );
  DFF_X1 reg_mem_reg_77__4_ ( .D(n6484), .CK(clk), .Q(n[1989]), .QN(n668) );
  DFF_X1 reg_mem_reg_77__3_ ( .D(n6483), .CK(clk), .Q(n[1988]), .QN(n669) );
  DFF_X1 reg_mem_reg_77__2_ ( .D(n6482), .CK(clk), .Q(n[1987]), .QN(n670) );
  DFF_X1 reg_mem_reg_77__1_ ( .D(n6481), .CK(clk), .Q(n[1986]), .QN(n671) );
  DFF_X1 reg_mem_reg_77__0_ ( .D(n6480), .CK(clk), .Q(n[1985]), .QN(n672) );
  DFF_X1 reg_mem_reg_78__7_ ( .D(n6479), .CK(clk), .QN(n689) );
  DFF_X1 reg_mem_reg_78__6_ ( .D(n6478), .CK(clk), .QN(n690) );
  DFF_X1 reg_mem_reg_78__5_ ( .D(n6477), .CK(clk), .QN(n691) );
  DFF_X1 reg_mem_reg_78__4_ ( .D(n6476), .CK(clk), .QN(n692) );
  DFF_X1 reg_mem_reg_78__3_ ( .D(n6475), .CK(clk), .QN(n693) );
  DFF_X1 reg_mem_reg_78__2_ ( .D(n6474), .CK(clk), .QN(n694) );
  DFF_X1 reg_mem_reg_78__1_ ( .D(n6473), .CK(clk), .QN(n695) );
  DFF_X1 reg_mem_reg_78__0_ ( .D(n6472), .CK(clk), .QN(n696) );
  DFF_X1 reg_mem_reg_79__7_ ( .D(n6471), .CK(clk), .QN(n697) );
  DFF_X1 reg_mem_reg_79__6_ ( .D(n6470), .CK(clk), .QN(n698) );
  DFF_X1 reg_mem_reg_79__5_ ( .D(n6469), .CK(clk), .QN(n699) );
  DFF_X1 reg_mem_reg_79__4_ ( .D(n6468), .CK(clk), .QN(n700) );
  DFF_X1 reg_mem_reg_79__3_ ( .D(n6467), .CK(clk), .QN(n701) );
  DFF_X1 reg_mem_reg_79__2_ ( .D(n6466), .CK(clk), .QN(n702) );
  DFF_X1 reg_mem_reg_79__1_ ( .D(n6465), .CK(clk), .QN(n703) );
  DFF_X1 reg_mem_reg_79__0_ ( .D(n6464), .CK(clk), .QN(n704) );
  DFF_X1 reg_mem_reg_80__7_ ( .D(n6463), .CK(clk), .Q(n[1968]), .QN(n721) );
  DFF_X1 reg_mem_reg_80__6_ ( .D(n6462), .CK(clk), .Q(n[1967]), .QN(n722) );
  DFF_X1 reg_mem_reg_80__5_ ( .D(n6461), .CK(clk), .Q(n[1966]), .QN(n723) );
  DFF_X1 reg_mem_reg_80__4_ ( .D(n6460), .CK(clk), .Q(n[1965]), .QN(n724) );
  DFF_X1 reg_mem_reg_80__3_ ( .D(n6459), .CK(clk), .Q(n[1964]), .QN(n725) );
  DFF_X1 reg_mem_reg_80__2_ ( .D(n6458), .CK(clk), .Q(n[1963]), .QN(n726) );
  DFF_X1 reg_mem_reg_80__1_ ( .D(n6457), .CK(clk), .Q(n[1962]), .QN(n727) );
  DFF_X1 reg_mem_reg_80__0_ ( .D(n6456), .CK(clk), .Q(n[1961]), .QN(n728) );
  DFF_X1 reg_mem_reg_81__7_ ( .D(n6455), .CK(clk), .Q(n[1960]), .QN(n729) );
  DFF_X1 reg_mem_reg_81__6_ ( .D(n6454), .CK(clk), .Q(n[1959]), .QN(n730) );
  DFF_X1 reg_mem_reg_81__5_ ( .D(n6453), .CK(clk), .Q(n[1958]), .QN(n731) );
  DFF_X1 reg_mem_reg_81__4_ ( .D(n6452), .CK(clk), .Q(n[1957]), .QN(n732) );
  DFF_X1 reg_mem_reg_81__3_ ( .D(n6451), .CK(clk), .Q(n[1956]), .QN(n733) );
  DFF_X1 reg_mem_reg_81__2_ ( .D(n6450), .CK(clk), .Q(n[1955]), .QN(n734) );
  DFF_X1 reg_mem_reg_81__1_ ( .D(n6449), .CK(clk), .Q(n[1954]), .QN(n735) );
  DFF_X1 reg_mem_reg_81__0_ ( .D(n6448), .CK(clk), .Q(n[1953]), .QN(n736) );
  DFF_X1 reg_mem_reg_82__7_ ( .D(n6447), .CK(clk), .QN(n753) );
  DFF_X1 reg_mem_reg_82__6_ ( .D(n6446), .CK(clk), .QN(n754) );
  DFF_X1 reg_mem_reg_82__5_ ( .D(n6445), .CK(clk), .QN(n755) );
  DFF_X1 reg_mem_reg_82__4_ ( .D(n6444), .CK(clk), .QN(n756) );
  DFF_X1 reg_mem_reg_82__3_ ( .D(n6443), .CK(clk), .QN(n757) );
  DFF_X1 reg_mem_reg_82__2_ ( .D(n6442), .CK(clk), .QN(n758) );
  DFF_X1 reg_mem_reg_82__1_ ( .D(n6441), .CK(clk), .QN(n759) );
  DFF_X1 reg_mem_reg_82__0_ ( .D(n6440), .CK(clk), .QN(n760) );
  DFF_X1 reg_mem_reg_83__7_ ( .D(n6439), .CK(clk), .QN(n761) );
  DFF_X1 reg_mem_reg_83__6_ ( .D(n6438), .CK(clk), .QN(n762) );
  DFF_X1 reg_mem_reg_83__5_ ( .D(n6437), .CK(clk), .QN(n763) );
  DFF_X1 reg_mem_reg_83__4_ ( .D(n6436), .CK(clk), .QN(n764) );
  DFF_X1 reg_mem_reg_83__3_ ( .D(n6435), .CK(clk), .QN(n765) );
  DFF_X1 reg_mem_reg_83__2_ ( .D(n6434), .CK(clk), .QN(n766) );
  DFF_X1 reg_mem_reg_83__1_ ( .D(n6433), .CK(clk), .QN(n767) );
  DFF_X1 reg_mem_reg_83__0_ ( .D(n6432), .CK(clk), .QN(n768) );
  DFF_X1 reg_mem_reg_84__7_ ( .D(n6431), .CK(clk), .Q(n[1936]), .QN(n785) );
  DFF_X1 reg_mem_reg_84__6_ ( .D(n6430), .CK(clk), .Q(n[1935]), .QN(n786) );
  DFF_X1 reg_mem_reg_84__5_ ( .D(n6429), .CK(clk), .Q(n[1934]), .QN(n787) );
  DFF_X1 reg_mem_reg_84__4_ ( .D(n6428), .CK(clk), .Q(n[1933]), .QN(n788) );
  DFF_X1 reg_mem_reg_84__3_ ( .D(n6427), .CK(clk), .Q(n[1932]), .QN(n789) );
  DFF_X1 reg_mem_reg_84__2_ ( .D(n6426), .CK(clk), .Q(n[1931]), .QN(n790) );
  DFF_X1 reg_mem_reg_84__1_ ( .D(n6425), .CK(clk), .Q(n[1930]), .QN(n791) );
  DFF_X1 reg_mem_reg_84__0_ ( .D(n6424), .CK(clk), .Q(n[1929]), .QN(n792) );
  DFF_X1 reg_mem_reg_85__7_ ( .D(n6423), .CK(clk), .Q(n[1928]), .QN(n793) );
  DFF_X1 reg_mem_reg_85__6_ ( .D(n6422), .CK(clk), .Q(n[1927]), .QN(n794) );
  DFF_X1 reg_mem_reg_85__5_ ( .D(n6421), .CK(clk), .Q(n[1926]), .QN(n795) );
  DFF_X1 reg_mem_reg_85__4_ ( .D(n6420), .CK(clk), .Q(n[1925]), .QN(n796) );
  DFF_X1 reg_mem_reg_85__3_ ( .D(n6419), .CK(clk), .Q(n[1924]), .QN(n797) );
  DFF_X1 reg_mem_reg_85__2_ ( .D(n6418), .CK(clk), .Q(n[1923]), .QN(n798) );
  DFF_X1 reg_mem_reg_85__1_ ( .D(n6417), .CK(clk), .Q(n[1922]), .QN(n799) );
  DFF_X1 reg_mem_reg_85__0_ ( .D(n6416), .CK(clk), .Q(n[1921]), .QN(n800) );
  DFF_X1 reg_mem_reg_86__7_ ( .D(n6415), .CK(clk), .QN(n817) );
  DFF_X1 reg_mem_reg_86__6_ ( .D(n6414), .CK(clk), .QN(n818) );
  DFF_X1 reg_mem_reg_86__5_ ( .D(n6413), .CK(clk), .QN(n819) );
  DFF_X1 reg_mem_reg_86__4_ ( .D(n6412), .CK(clk), .QN(n820) );
  DFF_X1 reg_mem_reg_86__3_ ( .D(n6411), .CK(clk), .QN(n821) );
  DFF_X1 reg_mem_reg_86__2_ ( .D(n6410), .CK(clk), .QN(n822) );
  DFF_X1 reg_mem_reg_86__1_ ( .D(n6409), .CK(clk), .QN(n823) );
  DFF_X1 reg_mem_reg_86__0_ ( .D(n6408), .CK(clk), .QN(n824) );
  DFF_X1 reg_mem_reg_87__7_ ( .D(n6407), .CK(clk), .QN(n825) );
  DFF_X1 reg_mem_reg_87__6_ ( .D(n6406), .CK(clk), .QN(n826) );
  DFF_X1 reg_mem_reg_87__5_ ( .D(n6405), .CK(clk), .QN(n827) );
  DFF_X1 reg_mem_reg_87__4_ ( .D(n6404), .CK(clk), .QN(n828) );
  DFF_X1 reg_mem_reg_87__3_ ( .D(n6403), .CK(clk), .QN(n829) );
  DFF_X1 reg_mem_reg_87__2_ ( .D(n6402), .CK(clk), .QN(n830) );
  DFF_X1 reg_mem_reg_87__1_ ( .D(n6401), .CK(clk), .QN(n831) );
  DFF_X1 reg_mem_reg_87__0_ ( .D(n6400), .CK(clk), .QN(n832) );
  DFF_X1 reg_mem_reg_88__7_ ( .D(n6399), .CK(clk), .Q(n[1904]), .QN(n849) );
  DFF_X1 reg_mem_reg_88__6_ ( .D(n6398), .CK(clk), .Q(n[1903]), .QN(n850) );
  DFF_X1 reg_mem_reg_88__5_ ( .D(n6397), .CK(clk), .Q(n[1902]), .QN(n851) );
  DFF_X1 reg_mem_reg_88__4_ ( .D(n6396), .CK(clk), .Q(n[1901]), .QN(n852) );
  DFF_X1 reg_mem_reg_88__3_ ( .D(n6395), .CK(clk), .Q(n[1900]), .QN(n853) );
  DFF_X1 reg_mem_reg_88__2_ ( .D(n6394), .CK(clk), .Q(n[1899]), .QN(n854) );
  DFF_X1 reg_mem_reg_88__1_ ( .D(n6393), .CK(clk), .Q(n[1898]), .QN(n855) );
  DFF_X1 reg_mem_reg_88__0_ ( .D(n6392), .CK(clk), .Q(n[1897]), .QN(n856) );
  DFF_X1 reg_mem_reg_89__7_ ( .D(n6391), .CK(clk), .Q(n[1896]), .QN(n857) );
  DFF_X1 reg_mem_reg_89__6_ ( .D(n6390), .CK(clk), .Q(n[1895]), .QN(n858) );
  DFF_X1 reg_mem_reg_89__5_ ( .D(n6389), .CK(clk), .Q(n[1894]), .QN(n859) );
  DFF_X1 reg_mem_reg_89__4_ ( .D(n6388), .CK(clk), .Q(n[1893]), .QN(n860) );
  DFF_X1 reg_mem_reg_89__3_ ( .D(n6387), .CK(clk), .Q(n[1892]), .QN(n861) );
  DFF_X1 reg_mem_reg_89__2_ ( .D(n6386), .CK(clk), .Q(n[1891]), .QN(n862) );
  DFF_X1 reg_mem_reg_89__1_ ( .D(n6385), .CK(clk), .Q(n[1890]), .QN(n863) );
  DFF_X1 reg_mem_reg_89__0_ ( .D(n6384), .CK(clk), .Q(n[1889]), .QN(n864) );
  DFF_X1 reg_mem_reg_90__7_ ( .D(n6383), .CK(clk), .QN(n881) );
  DFF_X1 reg_mem_reg_90__6_ ( .D(n6382), .CK(clk), .QN(n882) );
  DFF_X1 reg_mem_reg_90__5_ ( .D(n6381), .CK(clk), .QN(n883) );
  DFF_X1 reg_mem_reg_90__4_ ( .D(n6380), .CK(clk), .QN(n884) );
  DFF_X1 reg_mem_reg_90__3_ ( .D(n6379), .CK(clk), .QN(n885) );
  DFF_X1 reg_mem_reg_90__2_ ( .D(n6378), .CK(clk), .QN(n886) );
  DFF_X1 reg_mem_reg_90__1_ ( .D(n6377), .CK(clk), .QN(n887) );
  DFF_X1 reg_mem_reg_90__0_ ( .D(n6376), .CK(clk), .QN(n888) );
  DFF_X1 reg_mem_reg_91__7_ ( .D(n6375), .CK(clk), .QN(n889) );
  DFF_X1 reg_mem_reg_91__6_ ( .D(n6374), .CK(clk), .QN(n890) );
  DFF_X1 reg_mem_reg_91__5_ ( .D(n6373), .CK(clk), .QN(n891) );
  DFF_X1 reg_mem_reg_91__4_ ( .D(n6372), .CK(clk), .QN(n892) );
  DFF_X1 reg_mem_reg_91__3_ ( .D(n6371), .CK(clk), .QN(n893) );
  DFF_X1 reg_mem_reg_91__2_ ( .D(n6370), .CK(clk), .QN(n894) );
  DFF_X1 reg_mem_reg_91__1_ ( .D(n6369), .CK(clk), .QN(n895) );
  DFF_X1 reg_mem_reg_91__0_ ( .D(n6368), .CK(clk), .QN(n896) );
  DFF_X1 reg_mem_reg_92__7_ ( .D(n6367), .CK(clk), .Q(n[1872]), .QN(n913) );
  DFF_X1 reg_mem_reg_92__6_ ( .D(n6366), .CK(clk), .Q(n[1871]), .QN(n914) );
  DFF_X1 reg_mem_reg_92__5_ ( .D(n6365), .CK(clk), .Q(n[1870]), .QN(n915) );
  DFF_X1 reg_mem_reg_92__4_ ( .D(n6364), .CK(clk), .Q(n[1869]), .QN(n916) );
  DFF_X1 reg_mem_reg_92__3_ ( .D(n6363), .CK(clk), .Q(n[1868]), .QN(n917) );
  DFF_X1 reg_mem_reg_92__2_ ( .D(n6362), .CK(clk), .Q(n[1867]), .QN(n918) );
  DFF_X1 reg_mem_reg_92__1_ ( .D(n6361), .CK(clk), .Q(n[1866]), .QN(n919) );
  DFF_X1 reg_mem_reg_92__0_ ( .D(n6360), .CK(clk), .Q(n[1865]), .QN(n920) );
  DFF_X1 reg_mem_reg_93__7_ ( .D(n6359), .CK(clk), .Q(n[1864]), .QN(n921) );
  DFF_X1 reg_mem_reg_93__6_ ( .D(n6358), .CK(clk), .Q(n[1863]), .QN(n922) );
  DFF_X1 reg_mem_reg_93__5_ ( .D(n6357), .CK(clk), .Q(n[1862]), .QN(n923) );
  DFF_X1 reg_mem_reg_93__4_ ( .D(n6356), .CK(clk), .Q(n[1861]), .QN(n924) );
  DFF_X1 reg_mem_reg_93__3_ ( .D(n6355), .CK(clk), .Q(n[1860]), .QN(n925) );
  DFF_X1 reg_mem_reg_93__2_ ( .D(n6354), .CK(clk), .Q(n[1859]), .QN(n926) );
  DFF_X1 reg_mem_reg_93__1_ ( .D(n6353), .CK(clk), .Q(n[1858]), .QN(n927) );
  DFF_X1 reg_mem_reg_93__0_ ( .D(n6352), .CK(clk), .Q(n[1857]), .QN(n928) );
  DFF_X1 reg_mem_reg_94__7_ ( .D(n6351), .CK(clk), .QN(n945) );
  DFF_X1 reg_mem_reg_94__6_ ( .D(n6350), .CK(clk), .QN(n946) );
  DFF_X1 reg_mem_reg_94__5_ ( .D(n6349), .CK(clk), .QN(n947) );
  DFF_X1 reg_mem_reg_94__4_ ( .D(n6348), .CK(clk), .QN(n948) );
  DFF_X1 reg_mem_reg_94__3_ ( .D(n6347), .CK(clk), .QN(n949) );
  DFF_X1 reg_mem_reg_94__2_ ( .D(n6346), .CK(clk), .QN(n950) );
  DFF_X1 reg_mem_reg_94__1_ ( .D(n6345), .CK(clk), .QN(n951) );
  DFF_X1 reg_mem_reg_94__0_ ( .D(n6344), .CK(clk), .QN(n952) );
  DFF_X1 reg_mem_reg_95__7_ ( .D(n6343), .CK(clk), .QN(n953) );
  DFF_X1 reg_mem_reg_95__6_ ( .D(n6342), .CK(clk), .QN(n954) );
  DFF_X1 reg_mem_reg_95__5_ ( .D(n6341), .CK(clk), .QN(n955) );
  DFF_X1 reg_mem_reg_95__4_ ( .D(n6340), .CK(clk), .QN(n956) );
  DFF_X1 reg_mem_reg_95__3_ ( .D(n6339), .CK(clk), .QN(n957) );
  DFF_X1 reg_mem_reg_95__2_ ( .D(n6338), .CK(clk), .QN(n958) );
  DFF_X1 reg_mem_reg_95__1_ ( .D(n6337), .CK(clk), .QN(n959) );
  DFF_X1 reg_mem_reg_95__0_ ( .D(n6336), .CK(clk), .QN(n960) );
  DFF_X1 reg_mem_reg_96__7_ ( .D(n6335), .CK(clk), .Q(n[1840]), .QN(n977) );
  DFF_X1 reg_mem_reg_96__6_ ( .D(n6334), .CK(clk), .Q(n[1839]), .QN(n978) );
  DFF_X1 reg_mem_reg_96__5_ ( .D(n6333), .CK(clk), .Q(n[1838]), .QN(n979) );
  DFF_X1 reg_mem_reg_96__4_ ( .D(n6332), .CK(clk), .Q(n[1837]), .QN(n980) );
  DFF_X1 reg_mem_reg_96__3_ ( .D(n6331), .CK(clk), .Q(n[1836]), .QN(n981) );
  DFF_X1 reg_mem_reg_96__2_ ( .D(n6330), .CK(clk), .Q(n[1835]), .QN(n982) );
  DFF_X1 reg_mem_reg_96__1_ ( .D(n6329), .CK(clk), .Q(n[1834]), .QN(n983) );
  DFF_X1 reg_mem_reg_96__0_ ( .D(n6328), .CK(clk), .Q(n[1833]), .QN(n984) );
  DFF_X1 reg_mem_reg_97__7_ ( .D(n6327), .CK(clk), .Q(n[1832]), .QN(n985) );
  DFF_X1 reg_mem_reg_97__6_ ( .D(n6326), .CK(clk), .Q(n[1831]), .QN(n986) );
  DFF_X1 reg_mem_reg_97__5_ ( .D(n6325), .CK(clk), .Q(n[1830]), .QN(n987) );
  DFF_X1 reg_mem_reg_97__4_ ( .D(n6324), .CK(clk), .Q(n[1829]), .QN(n988) );
  DFF_X1 reg_mem_reg_97__3_ ( .D(n6323), .CK(clk), .Q(n[1828]), .QN(n989) );
  DFF_X1 reg_mem_reg_97__2_ ( .D(n6322), .CK(clk), .Q(n[1827]), .QN(n990) );
  DFF_X1 reg_mem_reg_97__1_ ( .D(n6321), .CK(clk), .Q(n[1826]), .QN(n991) );
  DFF_X1 reg_mem_reg_97__0_ ( .D(n6320), .CK(clk), .Q(n[1825]), .QN(n992) );
  DFF_X1 reg_mem_reg_98__7_ ( .D(n6319), .CK(clk), .QN(n1009) );
  DFF_X1 reg_mem_reg_98__6_ ( .D(n6318), .CK(clk), .QN(n1010) );
  DFF_X1 reg_mem_reg_98__5_ ( .D(n6317), .CK(clk), .QN(n1011) );
  DFF_X1 reg_mem_reg_98__4_ ( .D(n6316), .CK(clk), .QN(n1012) );
  DFF_X1 reg_mem_reg_98__3_ ( .D(n6315), .CK(clk), .QN(n1013) );
  DFF_X1 reg_mem_reg_98__2_ ( .D(n6314), .CK(clk), .QN(n1014) );
  DFF_X1 reg_mem_reg_98__1_ ( .D(n6313), .CK(clk), .QN(n1015) );
  DFF_X1 reg_mem_reg_98__0_ ( .D(n6312), .CK(clk), .QN(n1016) );
  DFF_X1 reg_mem_reg_99__7_ ( .D(n6311), .CK(clk), .QN(n1017) );
  DFF_X1 reg_mem_reg_99__6_ ( .D(n6310), .CK(clk), .QN(n1018) );
  DFF_X1 reg_mem_reg_99__5_ ( .D(n6309), .CK(clk), .QN(n1019) );
  DFF_X1 reg_mem_reg_99__4_ ( .D(n6308), .CK(clk), .QN(n1020) );
  DFF_X1 reg_mem_reg_99__3_ ( .D(n6307), .CK(clk), .QN(n1021) );
  DFF_X1 reg_mem_reg_99__2_ ( .D(n6306), .CK(clk), .QN(n1022) );
  DFF_X1 reg_mem_reg_99__1_ ( .D(n6305), .CK(clk), .QN(n1023) );
  DFF_X1 reg_mem_reg_99__0_ ( .D(n6304), .CK(clk), .QN(n1024) );
  DFF_X1 reg_mem_reg_100__7_ ( .D(n6303), .CK(clk), .Q(n[1808]), .QN(n1041) );
  DFF_X1 reg_mem_reg_100__6_ ( .D(n6302), .CK(clk), .Q(n[1807]), .QN(n1042) );
  DFF_X1 reg_mem_reg_100__5_ ( .D(n6301), .CK(clk), .Q(n[1806]), .QN(n1043) );
  DFF_X1 reg_mem_reg_100__4_ ( .D(n6300), .CK(clk), .Q(n[1805]), .QN(n1044) );
  DFF_X1 reg_mem_reg_100__3_ ( .D(n6299), .CK(clk), .Q(n[1804]), .QN(n1045) );
  DFF_X1 reg_mem_reg_100__2_ ( .D(n6298), .CK(clk), .Q(n[1803]), .QN(n1046) );
  DFF_X1 reg_mem_reg_100__1_ ( .D(n6297), .CK(clk), .Q(n[1802]), .QN(n1047) );
  DFF_X1 reg_mem_reg_100__0_ ( .D(n6296), .CK(clk), .Q(n[1801]), .QN(n1048) );
  DFF_X1 reg_mem_reg_101__7_ ( .D(n6295), .CK(clk), .Q(n[1800]), .QN(n1049) );
  DFF_X1 reg_mem_reg_101__6_ ( .D(n6294), .CK(clk), .Q(n[1799]), .QN(n1050) );
  DFF_X1 reg_mem_reg_101__5_ ( .D(n6293), .CK(clk), .Q(n[1798]), .QN(n1051) );
  DFF_X1 reg_mem_reg_101__4_ ( .D(n6292), .CK(clk), .Q(n[1797]), .QN(n1052) );
  DFF_X1 reg_mem_reg_101__3_ ( .D(n6291), .CK(clk), .Q(n[1796]), .QN(n1053) );
  DFF_X1 reg_mem_reg_101__2_ ( .D(n6290), .CK(clk), .Q(n[1795]), .QN(n1054) );
  DFF_X1 reg_mem_reg_101__1_ ( .D(n6289), .CK(clk), .Q(n[1794]), .QN(n1055) );
  DFF_X1 reg_mem_reg_101__0_ ( .D(n6288), .CK(clk), .Q(n[1793]), .QN(n1056) );
  DFF_X1 reg_mem_reg_102__7_ ( .D(n6287), .CK(clk), .QN(n1073) );
  DFF_X1 reg_mem_reg_102__6_ ( .D(n6286), .CK(clk), .QN(n1074) );
  DFF_X1 reg_mem_reg_102__5_ ( .D(n6285), .CK(clk), .QN(n1075) );
  DFF_X1 reg_mem_reg_102__4_ ( .D(n6284), .CK(clk), .QN(n1076) );
  DFF_X1 reg_mem_reg_102__3_ ( .D(n6283), .CK(clk), .QN(n1077) );
  DFF_X1 reg_mem_reg_102__2_ ( .D(n6282), .CK(clk), .QN(n1078) );
  DFF_X1 reg_mem_reg_102__1_ ( .D(n6281), .CK(clk), .QN(n1079) );
  DFF_X1 reg_mem_reg_102__0_ ( .D(n6280), .CK(clk), .QN(n1080) );
  DFF_X1 reg_mem_reg_103__7_ ( .D(n6279), .CK(clk), .QN(n1081) );
  DFF_X1 reg_mem_reg_103__6_ ( .D(n6278), .CK(clk), .QN(n1082) );
  DFF_X1 reg_mem_reg_103__5_ ( .D(n6277), .CK(clk), .QN(n1083) );
  DFF_X1 reg_mem_reg_103__4_ ( .D(n6276), .CK(clk), .QN(n1084) );
  DFF_X1 reg_mem_reg_103__3_ ( .D(n6275), .CK(clk), .QN(n1085) );
  DFF_X1 reg_mem_reg_103__2_ ( .D(n6274), .CK(clk), .QN(n1086) );
  DFF_X1 reg_mem_reg_103__1_ ( .D(n6273), .CK(clk), .QN(n1087) );
  DFF_X1 reg_mem_reg_103__0_ ( .D(n6272), .CK(clk), .QN(n1088) );
  DFF_X1 reg_mem_reg_104__7_ ( .D(n6271), .CK(clk), .Q(n[1776]), .QN(n1105) );
  DFF_X1 reg_mem_reg_104__6_ ( .D(n6270), .CK(clk), .Q(n[1775]), .QN(n1106) );
  DFF_X1 reg_mem_reg_104__5_ ( .D(n6269), .CK(clk), .Q(n[1774]), .QN(n1107) );
  DFF_X1 reg_mem_reg_104__4_ ( .D(n6268), .CK(clk), .Q(n[1773]), .QN(n1108) );
  DFF_X1 reg_mem_reg_104__3_ ( .D(n6267), .CK(clk), .Q(n[1772]), .QN(n1109) );
  DFF_X1 reg_mem_reg_104__2_ ( .D(n6266), .CK(clk), .Q(n[1771]), .QN(n1110) );
  DFF_X1 reg_mem_reg_104__1_ ( .D(n6265), .CK(clk), .Q(n[1770]), .QN(n1111) );
  DFF_X1 reg_mem_reg_104__0_ ( .D(n6264), .CK(clk), .Q(n[1769]), .QN(n1112) );
  DFF_X1 reg_mem_reg_105__7_ ( .D(n6263), .CK(clk), .Q(n[1768]), .QN(n1113) );
  DFF_X1 reg_mem_reg_105__6_ ( .D(n6262), .CK(clk), .Q(n[1767]), .QN(n1114) );
  DFF_X1 reg_mem_reg_105__5_ ( .D(n6261), .CK(clk), .Q(n[1766]), .QN(n1115) );
  DFF_X1 reg_mem_reg_105__4_ ( .D(n6260), .CK(clk), .Q(n[1765]), .QN(n1116) );
  DFF_X1 reg_mem_reg_105__3_ ( .D(n6259), .CK(clk), .Q(n[1764]), .QN(n1117) );
  DFF_X1 reg_mem_reg_105__2_ ( .D(n6258), .CK(clk), .Q(n[1763]), .QN(n1118) );
  DFF_X1 reg_mem_reg_105__1_ ( .D(n6257), .CK(clk), .Q(n[1762]), .QN(n1119) );
  DFF_X1 reg_mem_reg_105__0_ ( .D(n6256), .CK(clk), .Q(n[1761]), .QN(n1120) );
  DFF_X1 reg_mem_reg_106__7_ ( .D(n6255), .CK(clk), .QN(n1137) );
  DFF_X1 reg_mem_reg_106__6_ ( .D(n6254), .CK(clk), .QN(n1138) );
  DFF_X1 reg_mem_reg_106__5_ ( .D(n6253), .CK(clk), .QN(n1139) );
  DFF_X1 reg_mem_reg_106__4_ ( .D(n6252), .CK(clk), .QN(n1140) );
  DFF_X1 reg_mem_reg_106__3_ ( .D(n6251), .CK(clk), .QN(n1141) );
  DFF_X1 reg_mem_reg_106__2_ ( .D(n6250), .CK(clk), .QN(n1142) );
  DFF_X1 reg_mem_reg_106__1_ ( .D(n6249), .CK(clk), .QN(n1143) );
  DFF_X1 reg_mem_reg_106__0_ ( .D(n6248), .CK(clk), .QN(n1144) );
  DFF_X1 reg_mem_reg_107__7_ ( .D(n6247), .CK(clk), .QN(n1145) );
  DFF_X1 reg_mem_reg_107__6_ ( .D(n6246), .CK(clk), .QN(n1146) );
  DFF_X1 reg_mem_reg_107__5_ ( .D(n6245), .CK(clk), .QN(n1147) );
  DFF_X1 reg_mem_reg_107__4_ ( .D(n6244), .CK(clk), .QN(n1148) );
  DFF_X1 reg_mem_reg_107__3_ ( .D(n6243), .CK(clk), .QN(n1149) );
  DFF_X1 reg_mem_reg_107__2_ ( .D(n6242), .CK(clk), .QN(n1150) );
  DFF_X1 reg_mem_reg_107__1_ ( .D(n6241), .CK(clk), .QN(n1151) );
  DFF_X1 reg_mem_reg_107__0_ ( .D(n6240), .CK(clk), .QN(n1152) );
  DFF_X1 reg_mem_reg_108__7_ ( .D(n6239), .CK(clk), .Q(n[1744]), .QN(n1169) );
  DFF_X1 reg_mem_reg_108__6_ ( .D(n6238), .CK(clk), .Q(n[1743]), .QN(n1170) );
  DFF_X1 reg_mem_reg_108__5_ ( .D(n6237), .CK(clk), .Q(n[1742]), .QN(n1171) );
  DFF_X1 reg_mem_reg_108__4_ ( .D(n6236), .CK(clk), .Q(n[1741]), .QN(n1172) );
  DFF_X1 reg_mem_reg_108__3_ ( .D(n6235), .CK(clk), .Q(n[1740]), .QN(n1173) );
  DFF_X1 reg_mem_reg_108__2_ ( .D(n6234), .CK(clk), .Q(n[1739]), .QN(n1174) );
  DFF_X1 reg_mem_reg_108__1_ ( .D(n6233), .CK(clk), .Q(n[1738]), .QN(n1175) );
  DFF_X1 reg_mem_reg_108__0_ ( .D(n6232), .CK(clk), .Q(n[1737]), .QN(n1176) );
  DFF_X1 reg_mem_reg_109__7_ ( .D(n6231), .CK(clk), .Q(n[1736]), .QN(n1177) );
  DFF_X1 reg_mem_reg_109__6_ ( .D(n6230), .CK(clk), .Q(n[1735]), .QN(n1178) );
  DFF_X1 reg_mem_reg_109__5_ ( .D(n6229), .CK(clk), .Q(n[1734]), .QN(n1179) );
  DFF_X1 reg_mem_reg_109__4_ ( .D(n6228), .CK(clk), .Q(n[1733]), .QN(n1180) );
  DFF_X1 reg_mem_reg_109__3_ ( .D(n6227), .CK(clk), .Q(n[1732]), .QN(n1181) );
  DFF_X1 reg_mem_reg_109__2_ ( .D(n6226), .CK(clk), .Q(n[1731]), .QN(n1182) );
  DFF_X1 reg_mem_reg_109__1_ ( .D(n6225), .CK(clk), .Q(n[1730]), .QN(n1183) );
  DFF_X1 reg_mem_reg_109__0_ ( .D(n6224), .CK(clk), .Q(n[1729]), .QN(n1184) );
  DFF_X1 reg_mem_reg_110__7_ ( .D(n6223), .CK(clk), .QN(n1201) );
  DFF_X1 reg_mem_reg_110__6_ ( .D(n6222), .CK(clk), .QN(n1202) );
  DFF_X1 reg_mem_reg_110__5_ ( .D(n6221), .CK(clk), .QN(n1203) );
  DFF_X1 reg_mem_reg_110__4_ ( .D(n6220), .CK(clk), .QN(n1204) );
  DFF_X1 reg_mem_reg_110__3_ ( .D(n6219), .CK(clk), .QN(n1205) );
  DFF_X1 reg_mem_reg_110__2_ ( .D(n6218), .CK(clk), .QN(n1206) );
  DFF_X1 reg_mem_reg_110__1_ ( .D(n6217), .CK(clk), .QN(n1207) );
  DFF_X1 reg_mem_reg_110__0_ ( .D(n6216), .CK(clk), .QN(n1208) );
  DFF_X1 reg_mem_reg_111__7_ ( .D(n6215), .CK(clk), .QN(n1209) );
  DFF_X1 reg_mem_reg_111__6_ ( .D(n6214), .CK(clk), .QN(n1210) );
  DFF_X1 reg_mem_reg_111__5_ ( .D(n6213), .CK(clk), .QN(n1211) );
  DFF_X1 reg_mem_reg_111__4_ ( .D(n6212), .CK(clk), .QN(n1212) );
  DFF_X1 reg_mem_reg_111__3_ ( .D(n6211), .CK(clk), .QN(n1213) );
  DFF_X1 reg_mem_reg_111__2_ ( .D(n6210), .CK(clk), .QN(n1214) );
  DFF_X1 reg_mem_reg_111__1_ ( .D(n6209), .CK(clk), .QN(n1215) );
  DFF_X1 reg_mem_reg_111__0_ ( .D(n6208), .CK(clk), .QN(n1216) );
  DFF_X1 reg_mem_reg_112__7_ ( .D(n6207), .CK(clk), .Q(n[1712]), .QN(n1233) );
  DFF_X1 reg_mem_reg_112__6_ ( .D(n6206), .CK(clk), .Q(n[1711]), .QN(n1234) );
  DFF_X1 reg_mem_reg_112__5_ ( .D(n6205), .CK(clk), .Q(n[1710]), .QN(n1235) );
  DFF_X1 reg_mem_reg_112__4_ ( .D(n6204), .CK(clk), .Q(n[1709]), .QN(n1236) );
  DFF_X1 reg_mem_reg_112__3_ ( .D(n6203), .CK(clk), .Q(n[1708]), .QN(n1237) );
  DFF_X1 reg_mem_reg_112__2_ ( .D(n6202), .CK(clk), .Q(n[1707]), .QN(n1238) );
  DFF_X1 reg_mem_reg_112__1_ ( .D(n6201), .CK(clk), .Q(n[1706]), .QN(n1239) );
  DFF_X1 reg_mem_reg_112__0_ ( .D(n6200), .CK(clk), .Q(n[1705]), .QN(n1240) );
  DFF_X1 reg_mem_reg_113__7_ ( .D(n6199), .CK(clk), .Q(n[1704]), .QN(n1241) );
  DFF_X1 reg_mem_reg_113__6_ ( .D(n6198), .CK(clk), .Q(n[1703]), .QN(n1242) );
  DFF_X1 reg_mem_reg_113__5_ ( .D(n6197), .CK(clk), .Q(n[1702]), .QN(n1243) );
  DFF_X1 reg_mem_reg_113__4_ ( .D(n6196), .CK(clk), .Q(n[1701]), .QN(n1244) );
  DFF_X1 reg_mem_reg_113__3_ ( .D(n6195), .CK(clk), .Q(n[1700]), .QN(n1245) );
  DFF_X1 reg_mem_reg_113__2_ ( .D(n6194), .CK(clk), .Q(n[1699]), .QN(n1246) );
  DFF_X1 reg_mem_reg_113__1_ ( .D(n6193), .CK(clk), .Q(n[1698]), .QN(n1247) );
  DFF_X1 reg_mem_reg_113__0_ ( .D(n6192), .CK(clk), .Q(n[1697]), .QN(n1248) );
  DFF_X1 reg_mem_reg_114__7_ ( .D(n6191), .CK(clk), .QN(n1265) );
  DFF_X1 reg_mem_reg_114__6_ ( .D(n6190), .CK(clk), .QN(n1266) );
  DFF_X1 reg_mem_reg_114__5_ ( .D(n6189), .CK(clk), .QN(n1267) );
  DFF_X1 reg_mem_reg_114__4_ ( .D(n6188), .CK(clk), .QN(n1268) );
  DFF_X1 reg_mem_reg_114__3_ ( .D(n6187), .CK(clk), .QN(n1269) );
  DFF_X1 reg_mem_reg_114__2_ ( .D(n6186), .CK(clk), .QN(n1270) );
  DFF_X1 reg_mem_reg_114__1_ ( .D(n6185), .CK(clk), .QN(n1271) );
  DFF_X1 reg_mem_reg_114__0_ ( .D(n6184), .CK(clk), .QN(n1272) );
  DFF_X1 reg_mem_reg_115__7_ ( .D(n6183), .CK(clk), .QN(n1273) );
  DFF_X1 reg_mem_reg_115__6_ ( .D(n6182), .CK(clk), .QN(n1274) );
  DFF_X1 reg_mem_reg_115__5_ ( .D(n6181), .CK(clk), .QN(n1275) );
  DFF_X1 reg_mem_reg_115__4_ ( .D(n6180), .CK(clk), .QN(n1276) );
  DFF_X1 reg_mem_reg_115__3_ ( .D(n6179), .CK(clk), .QN(n1277) );
  DFF_X1 reg_mem_reg_115__2_ ( .D(n6178), .CK(clk), .QN(n1278) );
  DFF_X1 reg_mem_reg_115__1_ ( .D(n6177), .CK(clk), .QN(n1279) );
  DFF_X1 reg_mem_reg_115__0_ ( .D(n6176), .CK(clk), .QN(n1280) );
  DFF_X1 reg_mem_reg_116__7_ ( .D(n6175), .CK(clk), .Q(n[1680]), .QN(n1297) );
  DFF_X1 reg_mem_reg_116__6_ ( .D(n6174), .CK(clk), .Q(n[1679]), .QN(n1298) );
  DFF_X1 reg_mem_reg_116__5_ ( .D(n6173), .CK(clk), .Q(n[1678]), .QN(n1299) );
  DFF_X1 reg_mem_reg_116__4_ ( .D(n6172), .CK(clk), .Q(n[1677]), .QN(n1300) );
  DFF_X1 reg_mem_reg_116__3_ ( .D(n6171), .CK(clk), .Q(n[1676]), .QN(n1301) );
  DFF_X1 reg_mem_reg_116__2_ ( .D(n6170), .CK(clk), .Q(n[1675]), .QN(n1302) );
  DFF_X1 reg_mem_reg_116__1_ ( .D(n6169), .CK(clk), .Q(n[1674]), .QN(n1303) );
  DFF_X1 reg_mem_reg_116__0_ ( .D(n6168), .CK(clk), .Q(n[1673]), .QN(n1304) );
  DFF_X1 reg_mem_reg_117__7_ ( .D(n6167), .CK(clk), .Q(n[1672]), .QN(n1305) );
  DFF_X1 reg_mem_reg_117__6_ ( .D(n6166), .CK(clk), .Q(n[1671]), .QN(n1306) );
  DFF_X1 reg_mem_reg_117__5_ ( .D(n6165), .CK(clk), .Q(n[1670]), .QN(n1307) );
  DFF_X1 reg_mem_reg_117__4_ ( .D(n6164), .CK(clk), .Q(n[1669]), .QN(n1308) );
  DFF_X1 reg_mem_reg_117__3_ ( .D(n6163), .CK(clk), .Q(n[1668]), .QN(n1309) );
  DFF_X1 reg_mem_reg_117__2_ ( .D(n6162), .CK(clk), .Q(n[1667]), .QN(n1310) );
  DFF_X1 reg_mem_reg_117__1_ ( .D(n6161), .CK(clk), .Q(n[1666]), .QN(n1311) );
  DFF_X1 reg_mem_reg_117__0_ ( .D(n6160), .CK(clk), .Q(n[1665]), .QN(n1312) );
  DFF_X1 reg_mem_reg_118__7_ ( .D(n6159), .CK(clk), .QN(n1329) );
  DFF_X1 reg_mem_reg_118__6_ ( .D(n6158), .CK(clk), .QN(n1330) );
  DFF_X1 reg_mem_reg_118__5_ ( .D(n6157), .CK(clk), .QN(n1331) );
  DFF_X1 reg_mem_reg_118__4_ ( .D(n6156), .CK(clk), .QN(n1332) );
  DFF_X1 reg_mem_reg_118__3_ ( .D(n6155), .CK(clk), .QN(n1333) );
  DFF_X1 reg_mem_reg_118__2_ ( .D(n6154), .CK(clk), .QN(n1334) );
  DFF_X1 reg_mem_reg_118__1_ ( .D(n6153), .CK(clk), .QN(n1335) );
  DFF_X1 reg_mem_reg_118__0_ ( .D(n6152), .CK(clk), .QN(n1336) );
  DFF_X1 reg_mem_reg_119__7_ ( .D(n6151), .CK(clk), .QN(n1337) );
  DFF_X1 reg_mem_reg_119__6_ ( .D(n6150), .CK(clk), .QN(n1338) );
  DFF_X1 reg_mem_reg_119__5_ ( .D(n6149), .CK(clk), .QN(n1339) );
  DFF_X1 reg_mem_reg_119__4_ ( .D(n6148), .CK(clk), .QN(n1340) );
  DFF_X1 reg_mem_reg_119__3_ ( .D(n6147), .CK(clk), .QN(n1341) );
  DFF_X1 reg_mem_reg_119__2_ ( .D(n6146), .CK(clk), .QN(n1342) );
  DFF_X1 reg_mem_reg_119__1_ ( .D(n6145), .CK(clk), .QN(n1343) );
  DFF_X1 reg_mem_reg_119__0_ ( .D(n6144), .CK(clk), .QN(n1344) );
  DFF_X1 reg_mem_reg_120__7_ ( .D(n6143), .CK(clk), .Q(n[1648]), .QN(n1361) );
  DFF_X1 reg_mem_reg_120__6_ ( .D(n6142), .CK(clk), .Q(n[1647]), .QN(n1362) );
  DFF_X1 reg_mem_reg_120__5_ ( .D(n6141), .CK(clk), .Q(n[1646]), .QN(n1363) );
  DFF_X1 reg_mem_reg_120__4_ ( .D(n6140), .CK(clk), .Q(n[1645]), .QN(n1364) );
  DFF_X1 reg_mem_reg_120__3_ ( .D(n6139), .CK(clk), .Q(n[1644]), .QN(n1365) );
  DFF_X1 reg_mem_reg_120__2_ ( .D(n6138), .CK(clk), .Q(n[1643]), .QN(n1366) );
  DFF_X1 reg_mem_reg_120__1_ ( .D(n6137), .CK(clk), .Q(n[1642]), .QN(n1367) );
  DFF_X1 reg_mem_reg_120__0_ ( .D(n6136), .CK(clk), .Q(n[1641]), .QN(n1368) );
  DFF_X1 reg_mem_reg_121__7_ ( .D(n6135), .CK(clk), .Q(n[1640]), .QN(n1369) );
  DFF_X1 reg_mem_reg_121__6_ ( .D(n6134), .CK(clk), .Q(n[1639]), .QN(n1370) );
  DFF_X1 reg_mem_reg_121__5_ ( .D(n6133), .CK(clk), .Q(n[1638]), .QN(n1371) );
  DFF_X1 reg_mem_reg_121__4_ ( .D(n6132), .CK(clk), .Q(n[1637]), .QN(n1372) );
  DFF_X1 reg_mem_reg_121__3_ ( .D(n6131), .CK(clk), .Q(n[1636]), .QN(n1373) );
  DFF_X1 reg_mem_reg_121__2_ ( .D(n6130), .CK(clk), .Q(n[1635]), .QN(n1374) );
  DFF_X1 reg_mem_reg_121__1_ ( .D(n6129), .CK(clk), .Q(n[1634]), .QN(n1375) );
  DFF_X1 reg_mem_reg_121__0_ ( .D(n6128), .CK(clk), .Q(n[1633]), .QN(n1376) );
  DFF_X1 reg_mem_reg_122__7_ ( .D(n6127), .CK(clk), .QN(n1393) );
  DFF_X1 reg_mem_reg_122__6_ ( .D(n6126), .CK(clk), .QN(n1394) );
  DFF_X1 reg_mem_reg_122__5_ ( .D(n6125), .CK(clk), .QN(n1395) );
  DFF_X1 reg_mem_reg_122__4_ ( .D(n6124), .CK(clk), .QN(n1396) );
  DFF_X1 reg_mem_reg_122__3_ ( .D(n6123), .CK(clk), .QN(n1397) );
  DFF_X1 reg_mem_reg_122__2_ ( .D(n6122), .CK(clk), .QN(n1398) );
  DFF_X1 reg_mem_reg_122__1_ ( .D(n6121), .CK(clk), .QN(n1399) );
  DFF_X1 reg_mem_reg_122__0_ ( .D(n6120), .CK(clk), .QN(n1400) );
  DFF_X1 reg_mem_reg_123__7_ ( .D(n6119), .CK(clk), .QN(n1401) );
  DFF_X1 reg_mem_reg_123__6_ ( .D(n6118), .CK(clk), .QN(n1402) );
  DFF_X1 reg_mem_reg_123__5_ ( .D(n6117), .CK(clk), .QN(n1403) );
  DFF_X1 reg_mem_reg_123__4_ ( .D(n6116), .CK(clk), .QN(n1404) );
  DFF_X1 reg_mem_reg_123__3_ ( .D(n6115), .CK(clk), .QN(n1405) );
  DFF_X1 reg_mem_reg_123__2_ ( .D(n6114), .CK(clk), .QN(n1406) );
  DFF_X1 reg_mem_reg_123__1_ ( .D(n6113), .CK(clk), .QN(n1407) );
  DFF_X1 reg_mem_reg_123__0_ ( .D(n6112), .CK(clk), .QN(n1408) );
  DFF_X1 reg_mem_reg_124__7_ ( .D(n6111), .CK(clk), .Q(n[1616]), .QN(n1425) );
  DFF_X1 reg_mem_reg_124__6_ ( .D(n6110), .CK(clk), .Q(n[1615]), .QN(n1426) );
  DFF_X1 reg_mem_reg_124__5_ ( .D(n6109), .CK(clk), .Q(n[1614]), .QN(n1427) );
  DFF_X1 reg_mem_reg_124__4_ ( .D(n6108), .CK(clk), .Q(n[1613]), .QN(n1428) );
  DFF_X1 reg_mem_reg_124__3_ ( .D(n6107), .CK(clk), .Q(n[1612]), .QN(n1429) );
  DFF_X1 reg_mem_reg_124__2_ ( .D(n6106), .CK(clk), .Q(n[1611]), .QN(n1430) );
  DFF_X1 reg_mem_reg_124__1_ ( .D(n6105), .CK(clk), .Q(n[1610]), .QN(n1431) );
  DFF_X1 reg_mem_reg_124__0_ ( .D(n6104), .CK(clk), .Q(n[1609]), .QN(n1432) );
  DFF_X1 reg_mem_reg_125__7_ ( .D(n6103), .CK(clk), .Q(n[1608]), .QN(n1433) );
  DFF_X1 reg_mem_reg_125__6_ ( .D(n6102), .CK(clk), .Q(n[1607]), .QN(n1434) );
  DFF_X1 reg_mem_reg_125__5_ ( .D(n6101), .CK(clk), .Q(n[1606]), .QN(n1435) );
  DFF_X1 reg_mem_reg_125__4_ ( .D(n6100), .CK(clk), .Q(n[1605]), .QN(n1436) );
  DFF_X1 reg_mem_reg_125__3_ ( .D(n6099), .CK(clk), .Q(n[1604]), .QN(n1437) );
  DFF_X1 reg_mem_reg_125__2_ ( .D(n6098), .CK(clk), .Q(n[1603]), .QN(n1438) );
  DFF_X1 reg_mem_reg_125__1_ ( .D(n6097), .CK(clk), .Q(n[1602]), .QN(n1439) );
  DFF_X1 reg_mem_reg_125__0_ ( .D(n6096), .CK(clk), .Q(n[1601]), .QN(n1440) );
  DFF_X1 reg_mem_reg_126__7_ ( .D(n6095), .CK(clk), .QN(n1457) );
  DFF_X1 reg_mem_reg_126__6_ ( .D(n6094), .CK(clk), .QN(n1458) );
  DFF_X1 reg_mem_reg_126__5_ ( .D(n6093), .CK(clk), .QN(n1459) );
  DFF_X1 reg_mem_reg_126__4_ ( .D(n6092), .CK(clk), .QN(n1460) );
  DFF_X1 reg_mem_reg_126__3_ ( .D(n6091), .CK(clk), .QN(n1461) );
  DFF_X1 reg_mem_reg_126__2_ ( .D(n6090), .CK(clk), .QN(n1462) );
  DFF_X1 reg_mem_reg_126__1_ ( .D(n6089), .CK(clk), .QN(n1463) );
  DFF_X1 reg_mem_reg_126__0_ ( .D(n6088), .CK(clk), .QN(n1464) );
  DFF_X1 reg_mem_reg_127__7_ ( .D(n6087), .CK(clk), .QN(n1465) );
  DFF_X1 reg_mem_reg_127__6_ ( .D(n6086), .CK(clk), .QN(n1466) );
  DFF_X1 reg_mem_reg_127__5_ ( .D(n6085), .CK(clk), .QN(n1467) );
  DFF_X1 reg_mem_reg_127__4_ ( .D(n6084), .CK(clk), .QN(n1468) );
  DFF_X1 reg_mem_reg_127__3_ ( .D(n6083), .CK(clk), .QN(n1469) );
  DFF_X1 reg_mem_reg_127__2_ ( .D(n6082), .CK(clk), .QN(n1470) );
  DFF_X1 reg_mem_reg_127__1_ ( .D(n6081), .CK(clk), .QN(n1471) );
  DFF_X1 reg_mem_reg_127__0_ ( .D(n6080), .CK(clk), .QN(n1472) );
  DFF_X1 reg_mem_reg_128__7_ ( .D(n6079), .CK(clk), .Q(n[1584]), .QN(n1489) );
  DFF_X1 reg_mem_reg_128__6_ ( .D(n6078), .CK(clk), .Q(n[1583]), .QN(n1490) );
  DFF_X1 reg_mem_reg_128__5_ ( .D(n6077), .CK(clk), .Q(n[1582]), .QN(n1491) );
  DFF_X1 reg_mem_reg_128__4_ ( .D(n6076), .CK(clk), .Q(n[1581]), .QN(n1492) );
  DFF_X1 reg_mem_reg_128__3_ ( .D(n6075), .CK(clk), .Q(n[1580]), .QN(n1493) );
  DFF_X1 reg_mem_reg_128__2_ ( .D(n6074), .CK(clk), .Q(n[1579]), .QN(n1494) );
  DFF_X1 reg_mem_reg_128__1_ ( .D(n6073), .CK(clk), .Q(n[1578]), .QN(n1495) );
  DFF_X1 reg_mem_reg_128__0_ ( .D(n6072), .CK(clk), .Q(n[1577]), .QN(n1496) );
  DFF_X1 reg_mem_reg_129__7_ ( .D(n6071), .CK(clk), .Q(n[1576]), .QN(n1497) );
  DFF_X1 reg_mem_reg_129__6_ ( .D(n6070), .CK(clk), .Q(n[1575]), .QN(n1498) );
  DFF_X1 reg_mem_reg_129__5_ ( .D(n6069), .CK(clk), .Q(n[1574]), .QN(n1499) );
  DFF_X1 reg_mem_reg_129__4_ ( .D(n6068), .CK(clk), .Q(n[1573]), .QN(n1500) );
  DFF_X1 reg_mem_reg_129__3_ ( .D(n6067), .CK(clk), .Q(n[1572]), .QN(n1501) );
  DFF_X1 reg_mem_reg_129__2_ ( .D(n6066), .CK(clk), .Q(n[1571]), .QN(n1502) );
  DFF_X1 reg_mem_reg_129__1_ ( .D(n6065), .CK(clk), .Q(n[1570]), .QN(n1503) );
  DFF_X1 reg_mem_reg_129__0_ ( .D(n6064), .CK(clk), .Q(n[1569]), .QN(n1504) );
  DFF_X1 reg_mem_reg_130__7_ ( .D(n6063), .CK(clk), .QN(n1521) );
  DFF_X1 reg_mem_reg_130__6_ ( .D(n6062), .CK(clk), .QN(n1522) );
  DFF_X1 reg_mem_reg_130__5_ ( .D(n6061), .CK(clk), .QN(n1523) );
  DFF_X1 reg_mem_reg_130__4_ ( .D(n6060), .CK(clk), .QN(n1524) );
  DFF_X1 reg_mem_reg_130__3_ ( .D(n6059), .CK(clk), .QN(n1525) );
  DFF_X1 reg_mem_reg_130__2_ ( .D(n6058), .CK(clk), .QN(n1526) );
  DFF_X1 reg_mem_reg_130__1_ ( .D(n6057), .CK(clk), .QN(n1527) );
  DFF_X1 reg_mem_reg_130__0_ ( .D(n6056), .CK(clk), .QN(n1528) );
  DFF_X1 reg_mem_reg_131__7_ ( .D(n6055), .CK(clk), .QN(n1529) );
  DFF_X1 reg_mem_reg_131__6_ ( .D(n6054), .CK(clk), .QN(n1530) );
  DFF_X1 reg_mem_reg_131__5_ ( .D(n6053), .CK(clk), .QN(n1531) );
  DFF_X1 reg_mem_reg_131__4_ ( .D(n6052), .CK(clk), .QN(n1532) );
  DFF_X1 reg_mem_reg_131__3_ ( .D(n6051), .CK(clk), .QN(n1533) );
  DFF_X1 reg_mem_reg_131__2_ ( .D(n6050), .CK(clk), .QN(n1534) );
  DFF_X1 reg_mem_reg_131__1_ ( .D(n6049), .CK(clk), .QN(n1535) );
  DFF_X1 reg_mem_reg_131__0_ ( .D(n6048), .CK(clk), .QN(n1536) );
  DFF_X1 reg_mem_reg_132__7_ ( .D(n6047), .CK(clk), .Q(n[1552]), .QN(n1553) );
  DFF_X1 reg_mem_reg_132__6_ ( .D(n6046), .CK(clk), .Q(n[1551]), .QN(n1554) );
  DFF_X1 reg_mem_reg_132__5_ ( .D(n6045), .CK(clk), .Q(n[1550]), .QN(n1555) );
  DFF_X1 reg_mem_reg_132__4_ ( .D(n6044), .CK(clk), .Q(n[1549]), .QN(n1556) );
  DFF_X1 reg_mem_reg_132__3_ ( .D(n6043), .CK(clk), .Q(n[1548]), .QN(n1557) );
  DFF_X1 reg_mem_reg_132__2_ ( .D(n6042), .CK(clk), .Q(n[1547]), .QN(n1558) );
  DFF_X1 reg_mem_reg_132__1_ ( .D(n6041), .CK(clk), .Q(n[1546]), .QN(n1559) );
  DFF_X1 reg_mem_reg_132__0_ ( .D(n6040), .CK(clk), .Q(n[1545]), .QN(n1560) );
  DFF_X1 reg_mem_reg_133__7_ ( .D(n6039), .CK(clk), .Q(n[1544]), .QN(n1561) );
  DFF_X1 reg_mem_reg_133__6_ ( .D(n6038), .CK(clk), .Q(n[1543]), .QN(n1562) );
  DFF_X1 reg_mem_reg_133__5_ ( .D(n6037), .CK(clk), .Q(n[1542]), .QN(n1563) );
  DFF_X1 reg_mem_reg_133__4_ ( .D(n6036), .CK(clk), .Q(n[1541]), .QN(n1564) );
  DFF_X1 reg_mem_reg_133__3_ ( .D(n6035), .CK(clk), .Q(n[1540]), .QN(n1565) );
  DFF_X1 reg_mem_reg_133__2_ ( .D(n6034), .CK(clk), .Q(n[1539]), .QN(n1566) );
  DFF_X1 reg_mem_reg_133__1_ ( .D(n6033), .CK(clk), .Q(n[1538]), .QN(n1567) );
  DFF_X1 reg_mem_reg_133__0_ ( .D(n6032), .CK(clk), .Q(n[1537]), .QN(n1568) );
  DFF_X1 reg_mem_reg_134__7_ ( .D(n6031), .CK(clk), .QN(n1585) );
  DFF_X1 reg_mem_reg_134__6_ ( .D(n6030), .CK(clk), .QN(n1586) );
  DFF_X1 reg_mem_reg_134__5_ ( .D(n6029), .CK(clk), .QN(n1587) );
  DFF_X1 reg_mem_reg_134__4_ ( .D(n6028), .CK(clk), .QN(n1588) );
  DFF_X1 reg_mem_reg_134__3_ ( .D(n6027), .CK(clk), .QN(n1589) );
  DFF_X1 reg_mem_reg_134__2_ ( .D(n6026), .CK(clk), .QN(n1590) );
  DFF_X1 reg_mem_reg_134__1_ ( .D(n6025), .CK(clk), .QN(n1591) );
  DFF_X1 reg_mem_reg_134__0_ ( .D(n6024), .CK(clk), .QN(n1592) );
  DFF_X1 reg_mem_reg_135__7_ ( .D(n6023), .CK(clk), .QN(n1593) );
  DFF_X1 reg_mem_reg_135__6_ ( .D(n6022), .CK(clk), .QN(n1594) );
  DFF_X1 reg_mem_reg_135__5_ ( .D(n6021), .CK(clk), .QN(n1595) );
  DFF_X1 reg_mem_reg_135__4_ ( .D(n6020), .CK(clk), .QN(n1596) );
  DFF_X1 reg_mem_reg_135__3_ ( .D(n6019), .CK(clk), .QN(n1597) );
  DFF_X1 reg_mem_reg_135__2_ ( .D(n6018), .CK(clk), .QN(n1598) );
  DFF_X1 reg_mem_reg_135__1_ ( .D(n6017), .CK(clk), .QN(n1599) );
  DFF_X1 reg_mem_reg_135__0_ ( .D(n6016), .CK(clk), .QN(n1600) );
  DFF_X1 reg_mem_reg_136__7_ ( .D(n6015), .CK(clk), .Q(n[1520]), .QN(n1617) );
  DFF_X1 reg_mem_reg_136__6_ ( .D(n6014), .CK(clk), .Q(n[1519]), .QN(n1618) );
  DFF_X1 reg_mem_reg_136__5_ ( .D(n6013), .CK(clk), .Q(n[1518]), .QN(n1619) );
  DFF_X1 reg_mem_reg_136__4_ ( .D(n6012), .CK(clk), .Q(n[1517]), .QN(n1620) );
  DFF_X1 reg_mem_reg_136__3_ ( .D(n6011), .CK(clk), .Q(n[1516]), .QN(n1621) );
  DFF_X1 reg_mem_reg_136__2_ ( .D(n6010), .CK(clk), .Q(n[1515]), .QN(n1622) );
  DFF_X1 reg_mem_reg_136__1_ ( .D(n6009), .CK(clk), .Q(n[1514]), .QN(n1623) );
  DFF_X1 reg_mem_reg_136__0_ ( .D(n6008), .CK(clk), .Q(n[1513]), .QN(n1624) );
  DFF_X1 reg_mem_reg_137__7_ ( .D(n6007), .CK(clk), .Q(n[1512]), .QN(n1625) );
  DFF_X1 reg_mem_reg_137__6_ ( .D(n6006), .CK(clk), .Q(n[1511]), .QN(n1626) );
  DFF_X1 reg_mem_reg_137__5_ ( .D(n6005), .CK(clk), .Q(n[1510]), .QN(n1627) );
  DFF_X1 reg_mem_reg_137__4_ ( .D(n6004), .CK(clk), .Q(n[1509]), .QN(n1628) );
  DFF_X1 reg_mem_reg_137__3_ ( .D(n6003), .CK(clk), .Q(n[1508]), .QN(n1629) );
  DFF_X1 reg_mem_reg_137__2_ ( .D(n6002), .CK(clk), .Q(n[1507]), .QN(n1630) );
  DFF_X1 reg_mem_reg_137__1_ ( .D(n6001), .CK(clk), .Q(n[1506]), .QN(n1631) );
  DFF_X1 reg_mem_reg_137__0_ ( .D(n6000), .CK(clk), .Q(n[1505]), .QN(n1632) );
  DFF_X1 reg_mem_reg_138__7_ ( .D(n5999), .CK(clk), .QN(n1649) );
  DFF_X1 reg_mem_reg_138__6_ ( .D(n5998), .CK(clk), .QN(n1650) );
  DFF_X1 reg_mem_reg_138__5_ ( .D(n5997), .CK(clk), .QN(n1651) );
  DFF_X1 reg_mem_reg_138__4_ ( .D(n5996), .CK(clk), .QN(n1652) );
  DFF_X1 reg_mem_reg_138__3_ ( .D(n5995), .CK(clk), .QN(n1653) );
  DFF_X1 reg_mem_reg_138__2_ ( .D(n5994), .CK(clk), .QN(n1654) );
  DFF_X1 reg_mem_reg_138__1_ ( .D(n5993), .CK(clk), .QN(n1655) );
  DFF_X1 reg_mem_reg_138__0_ ( .D(n5992), .CK(clk), .QN(n1656) );
  DFF_X1 reg_mem_reg_139__7_ ( .D(n5991), .CK(clk), .QN(n1657) );
  DFF_X1 reg_mem_reg_139__6_ ( .D(n5990), .CK(clk), .QN(n1658) );
  DFF_X1 reg_mem_reg_139__5_ ( .D(n5989), .CK(clk), .QN(n1659) );
  DFF_X1 reg_mem_reg_139__4_ ( .D(n5988), .CK(clk), .QN(n1660) );
  DFF_X1 reg_mem_reg_139__3_ ( .D(n5987), .CK(clk), .QN(n1661) );
  DFF_X1 reg_mem_reg_139__2_ ( .D(n5986), .CK(clk), .QN(n1662) );
  DFF_X1 reg_mem_reg_139__1_ ( .D(n5985), .CK(clk), .QN(n1663) );
  DFF_X1 reg_mem_reg_139__0_ ( .D(n5984), .CK(clk), .QN(n1664) );
  DFF_X1 reg_mem_reg_140__7_ ( .D(n5983), .CK(clk), .Q(n[1488]), .QN(n1681) );
  DFF_X1 reg_mem_reg_140__6_ ( .D(n5982), .CK(clk), .Q(n[1487]), .QN(n1682) );
  DFF_X1 reg_mem_reg_140__5_ ( .D(n5981), .CK(clk), .Q(n[1486]), .QN(n1683) );
  DFF_X1 reg_mem_reg_140__4_ ( .D(n5980), .CK(clk), .Q(n[1485]), .QN(n1684) );
  DFF_X1 reg_mem_reg_140__3_ ( .D(n5979), .CK(clk), .Q(n[1484]), .QN(n1685) );
  DFF_X1 reg_mem_reg_140__2_ ( .D(n5978), .CK(clk), .Q(n[1483]), .QN(n1686) );
  DFF_X1 reg_mem_reg_140__1_ ( .D(n5977), .CK(clk), .Q(n[1482]), .QN(n1687) );
  DFF_X1 reg_mem_reg_140__0_ ( .D(n5976), .CK(clk), .Q(n[1481]), .QN(n1688) );
  DFF_X1 reg_mem_reg_141__7_ ( .D(n5975), .CK(clk), .Q(n[1480]), .QN(n1689) );
  DFF_X1 reg_mem_reg_141__6_ ( .D(n5974), .CK(clk), .Q(n[1479]), .QN(n1690) );
  DFF_X1 reg_mem_reg_141__5_ ( .D(n5973), .CK(clk), .Q(n[1478]), .QN(n1691) );
  DFF_X1 reg_mem_reg_141__4_ ( .D(n5972), .CK(clk), .Q(n[1477]), .QN(n1692) );
  DFF_X1 reg_mem_reg_141__3_ ( .D(n5971), .CK(clk), .Q(n[1476]), .QN(n1693) );
  DFF_X1 reg_mem_reg_141__2_ ( .D(n5970), .CK(clk), .Q(n[1475]), .QN(n1694) );
  DFF_X1 reg_mem_reg_141__1_ ( .D(n5969), .CK(clk), .Q(n[1474]), .QN(n1695) );
  DFF_X1 reg_mem_reg_141__0_ ( .D(n5968), .CK(clk), .Q(n[1473]), .QN(n1696) );
  DFF_X1 reg_mem_reg_142__7_ ( .D(n5967), .CK(clk), .QN(n1713) );
  DFF_X1 reg_mem_reg_142__6_ ( .D(n5966), .CK(clk), .QN(n1714) );
  DFF_X1 reg_mem_reg_142__5_ ( .D(n5965), .CK(clk), .QN(n1715) );
  DFF_X1 reg_mem_reg_142__4_ ( .D(n5964), .CK(clk), .QN(n1716) );
  DFF_X1 reg_mem_reg_142__3_ ( .D(n5963), .CK(clk), .QN(n1717) );
  DFF_X1 reg_mem_reg_142__2_ ( .D(n5962), .CK(clk), .QN(n1718) );
  DFF_X1 reg_mem_reg_142__1_ ( .D(n5961), .CK(clk), .QN(n1719) );
  DFF_X1 reg_mem_reg_142__0_ ( .D(n5960), .CK(clk), .QN(n1720) );
  DFF_X1 reg_mem_reg_143__7_ ( .D(n5959), .CK(clk), .QN(n1721) );
  DFF_X1 reg_mem_reg_143__6_ ( .D(n5958), .CK(clk), .QN(n1722) );
  DFF_X1 reg_mem_reg_143__5_ ( .D(n5957), .CK(clk), .QN(n1723) );
  DFF_X1 reg_mem_reg_143__4_ ( .D(n5956), .CK(clk), .QN(n1724) );
  DFF_X1 reg_mem_reg_143__3_ ( .D(n5955), .CK(clk), .QN(n1725) );
  DFF_X1 reg_mem_reg_143__2_ ( .D(n5954), .CK(clk), .QN(n1726) );
  DFF_X1 reg_mem_reg_143__1_ ( .D(n5953), .CK(clk), .QN(n1727) );
  DFF_X1 reg_mem_reg_143__0_ ( .D(n5952), .CK(clk), .QN(n1728) );
  DFF_X1 reg_mem_reg_144__7_ ( .D(n5951), .CK(clk), .Q(n[1456]), .QN(n1745) );
  DFF_X1 reg_mem_reg_144__6_ ( .D(n5950), .CK(clk), .Q(n[1455]), .QN(n1746) );
  DFF_X1 reg_mem_reg_144__5_ ( .D(n5949), .CK(clk), .Q(n[1454]), .QN(n1747) );
  DFF_X1 reg_mem_reg_144__4_ ( .D(n5948), .CK(clk), .Q(n[1453]), .QN(n1748) );
  DFF_X1 reg_mem_reg_144__3_ ( .D(n5947), .CK(clk), .Q(n[1452]), .QN(n1749) );
  DFF_X1 reg_mem_reg_144__2_ ( .D(n5946), .CK(clk), .Q(n[1451]), .QN(n1750) );
  DFF_X1 reg_mem_reg_144__1_ ( .D(n5945), .CK(clk), .Q(n[1450]), .QN(n1751) );
  DFF_X1 reg_mem_reg_144__0_ ( .D(n5944), .CK(clk), .Q(n[1449]), .QN(n1752) );
  DFF_X1 reg_mem_reg_145__7_ ( .D(n5943), .CK(clk), .Q(n[1448]), .QN(n1753) );
  DFF_X1 reg_mem_reg_145__6_ ( .D(n5942), .CK(clk), .Q(n[1447]), .QN(n1754) );
  DFF_X1 reg_mem_reg_145__5_ ( .D(n5941), .CK(clk), .Q(n[1446]), .QN(n1755) );
  DFF_X1 reg_mem_reg_145__4_ ( .D(n5940), .CK(clk), .Q(n[1445]), .QN(n1756) );
  DFF_X1 reg_mem_reg_145__3_ ( .D(n5939), .CK(clk), .Q(n[1444]), .QN(n1757) );
  DFF_X1 reg_mem_reg_145__2_ ( .D(n5938), .CK(clk), .Q(n[1443]), .QN(n1758) );
  DFF_X1 reg_mem_reg_145__1_ ( .D(n5937), .CK(clk), .Q(n[1442]), .QN(n1759) );
  DFF_X1 reg_mem_reg_145__0_ ( .D(n5936), .CK(clk), .Q(n[1441]), .QN(n1760) );
  DFF_X1 reg_mem_reg_146__7_ ( .D(n5935), .CK(clk), .QN(n1777) );
  DFF_X1 reg_mem_reg_146__6_ ( .D(n5934), .CK(clk), .QN(n1778) );
  DFF_X1 reg_mem_reg_146__5_ ( .D(n5933), .CK(clk), .QN(n1779) );
  DFF_X1 reg_mem_reg_146__4_ ( .D(n5932), .CK(clk), .QN(n1780) );
  DFF_X1 reg_mem_reg_146__3_ ( .D(n5931), .CK(clk), .QN(n1781) );
  DFF_X1 reg_mem_reg_146__2_ ( .D(n5930), .CK(clk), .QN(n1782) );
  DFF_X1 reg_mem_reg_146__1_ ( .D(n5929), .CK(clk), .QN(n1783) );
  DFF_X1 reg_mem_reg_146__0_ ( .D(n5928), .CK(clk), .QN(n1784) );
  DFF_X1 reg_mem_reg_147__7_ ( .D(n5927), .CK(clk), .QN(n1785) );
  DFF_X1 reg_mem_reg_147__6_ ( .D(n5926), .CK(clk), .QN(n1786) );
  DFF_X1 reg_mem_reg_147__5_ ( .D(n5925), .CK(clk), .QN(n1787) );
  DFF_X1 reg_mem_reg_147__4_ ( .D(n5924), .CK(clk), .QN(n1788) );
  DFF_X1 reg_mem_reg_147__3_ ( .D(n5923), .CK(clk), .QN(n1789) );
  DFF_X1 reg_mem_reg_147__2_ ( .D(n5922), .CK(clk), .QN(n1790) );
  DFF_X1 reg_mem_reg_147__1_ ( .D(n5921), .CK(clk), .QN(n1791) );
  DFF_X1 reg_mem_reg_147__0_ ( .D(n5920), .CK(clk), .QN(n1792) );
  DFF_X1 reg_mem_reg_148__7_ ( .D(n5919), .CK(clk), .Q(n[1424]), .QN(n1809) );
  DFF_X1 reg_mem_reg_148__6_ ( .D(n5918), .CK(clk), .Q(n[1423]), .QN(n1810) );
  DFF_X1 reg_mem_reg_148__5_ ( .D(n5917), .CK(clk), .Q(n[1422]), .QN(n1811) );
  DFF_X1 reg_mem_reg_148__4_ ( .D(n5916), .CK(clk), .Q(n[1421]), .QN(n1812) );
  DFF_X1 reg_mem_reg_148__3_ ( .D(n5915), .CK(clk), .Q(n[1420]), .QN(n1813) );
  DFF_X1 reg_mem_reg_148__2_ ( .D(n5914), .CK(clk), .Q(n[1419]), .QN(n1814) );
  DFF_X1 reg_mem_reg_148__1_ ( .D(n5913), .CK(clk), .Q(n[1418]), .QN(n1815) );
  DFF_X1 reg_mem_reg_148__0_ ( .D(n5912), .CK(clk), .Q(n[1417]), .QN(n1816) );
  DFF_X1 reg_mem_reg_149__7_ ( .D(n5911), .CK(clk), .Q(n[1416]), .QN(n1817) );
  DFF_X1 reg_mem_reg_149__6_ ( .D(n5910), .CK(clk), .Q(n[1415]), .QN(n1818) );
  DFF_X1 reg_mem_reg_149__5_ ( .D(n5909), .CK(clk), .Q(n[1414]), .QN(n1819) );
  DFF_X1 reg_mem_reg_149__4_ ( .D(n5908), .CK(clk), .Q(n[1413]), .QN(n1820) );
  DFF_X1 reg_mem_reg_149__3_ ( .D(n5907), .CK(clk), .Q(n[1412]), .QN(n1821) );
  DFF_X1 reg_mem_reg_149__2_ ( .D(n5906), .CK(clk), .Q(n[1411]), .QN(n1822) );
  DFF_X1 reg_mem_reg_149__1_ ( .D(n5905), .CK(clk), .Q(n[1410]), .QN(n1823) );
  DFF_X1 reg_mem_reg_149__0_ ( .D(n5904), .CK(clk), .Q(n[1409]), .QN(n1824) );
  DFF_X1 reg_mem_reg_150__7_ ( .D(n5903), .CK(clk), .QN(n1841) );
  DFF_X1 reg_mem_reg_150__6_ ( .D(n5902), .CK(clk), .QN(n1842) );
  DFF_X1 reg_mem_reg_150__5_ ( .D(n5901), .CK(clk), .QN(n1843) );
  DFF_X1 reg_mem_reg_150__4_ ( .D(n5900), .CK(clk), .QN(n1844) );
  DFF_X1 reg_mem_reg_150__3_ ( .D(n5899), .CK(clk), .QN(n1845) );
  DFF_X1 reg_mem_reg_150__2_ ( .D(n5898), .CK(clk), .QN(n1846) );
  DFF_X1 reg_mem_reg_150__1_ ( .D(n5897), .CK(clk), .QN(n1847) );
  DFF_X1 reg_mem_reg_150__0_ ( .D(n5896), .CK(clk), .QN(n1848) );
  DFF_X1 reg_mem_reg_151__7_ ( .D(n5895), .CK(clk), .QN(n1849) );
  DFF_X1 reg_mem_reg_151__6_ ( .D(n5894), .CK(clk), .QN(n1850) );
  DFF_X1 reg_mem_reg_151__5_ ( .D(n5893), .CK(clk), .QN(n1851) );
  DFF_X1 reg_mem_reg_151__4_ ( .D(n5892), .CK(clk), .QN(n1852) );
  DFF_X1 reg_mem_reg_151__3_ ( .D(n5891), .CK(clk), .QN(n1853) );
  DFF_X1 reg_mem_reg_151__2_ ( .D(n5890), .CK(clk), .QN(n1854) );
  DFF_X1 reg_mem_reg_151__1_ ( .D(n5889), .CK(clk), .QN(n1855) );
  DFF_X1 reg_mem_reg_151__0_ ( .D(n5888), .CK(clk), .QN(n1856) );
  DFF_X1 reg_mem_reg_152__7_ ( .D(n5887), .CK(clk), .Q(n[1392]), .QN(n1873) );
  DFF_X1 reg_mem_reg_152__6_ ( .D(n5886), .CK(clk), .Q(n[1391]), .QN(n1874) );
  DFF_X1 reg_mem_reg_152__5_ ( .D(n5885), .CK(clk), .Q(n[1390]), .QN(n1875) );
  DFF_X1 reg_mem_reg_152__4_ ( .D(n5884), .CK(clk), .Q(n[1389]), .QN(n1876) );
  DFF_X1 reg_mem_reg_152__3_ ( .D(n5883), .CK(clk), .Q(n[1388]), .QN(n1877) );
  DFF_X1 reg_mem_reg_152__2_ ( .D(n5882), .CK(clk), .Q(n[1387]), .QN(n1878) );
  DFF_X1 reg_mem_reg_152__1_ ( .D(n5881), .CK(clk), .Q(n[1386]), .QN(n1879) );
  DFF_X1 reg_mem_reg_152__0_ ( .D(n5880), .CK(clk), .Q(n[1385]), .QN(n1880) );
  DFF_X1 reg_mem_reg_153__7_ ( .D(n5879), .CK(clk), .Q(n[1384]), .QN(n1881) );
  DFF_X1 reg_mem_reg_153__6_ ( .D(n5878), .CK(clk), .Q(n[1383]), .QN(n1882) );
  DFF_X1 reg_mem_reg_153__5_ ( .D(n5877), .CK(clk), .Q(n[1382]), .QN(n1883) );
  DFF_X1 reg_mem_reg_153__4_ ( .D(n5876), .CK(clk), .Q(n[1381]), .QN(n1884) );
  DFF_X1 reg_mem_reg_153__3_ ( .D(n5875), .CK(clk), .Q(n[1380]), .QN(n1885) );
  DFF_X1 reg_mem_reg_153__2_ ( .D(n5874), .CK(clk), .Q(n[1379]), .QN(n1886) );
  DFF_X1 reg_mem_reg_153__1_ ( .D(n5873), .CK(clk), .Q(n[1378]), .QN(n1887) );
  DFF_X1 reg_mem_reg_153__0_ ( .D(n5872), .CK(clk), .Q(n[1377]), .QN(n1888) );
  DFF_X1 reg_mem_reg_154__7_ ( .D(n5871), .CK(clk), .QN(n1905) );
  DFF_X1 reg_mem_reg_154__6_ ( .D(n5870), .CK(clk), .QN(n1906) );
  DFF_X1 reg_mem_reg_154__5_ ( .D(n5869), .CK(clk), .QN(n1907) );
  DFF_X1 reg_mem_reg_154__4_ ( .D(n5868), .CK(clk), .QN(n1908) );
  DFF_X1 reg_mem_reg_154__3_ ( .D(n5867), .CK(clk), .QN(n1909) );
  DFF_X1 reg_mem_reg_154__2_ ( .D(n5866), .CK(clk), .QN(n1910) );
  DFF_X1 reg_mem_reg_154__1_ ( .D(n5865), .CK(clk), .QN(n1911) );
  DFF_X1 reg_mem_reg_154__0_ ( .D(n5864), .CK(clk), .QN(n1912) );
  DFF_X1 reg_mem_reg_155__7_ ( .D(n5863), .CK(clk), .QN(n1913) );
  DFF_X1 reg_mem_reg_155__6_ ( .D(n5862), .CK(clk), .QN(n1914) );
  DFF_X1 reg_mem_reg_155__5_ ( .D(n5861), .CK(clk), .QN(n1915) );
  DFF_X1 reg_mem_reg_155__4_ ( .D(n5860), .CK(clk), .QN(n1916) );
  DFF_X1 reg_mem_reg_155__3_ ( .D(n5859), .CK(clk), .QN(n1917) );
  DFF_X1 reg_mem_reg_155__2_ ( .D(n5858), .CK(clk), .QN(n1918) );
  DFF_X1 reg_mem_reg_155__1_ ( .D(n5857), .CK(clk), .QN(n1919) );
  DFF_X1 reg_mem_reg_155__0_ ( .D(n5856), .CK(clk), .QN(n1920) );
  DFF_X1 reg_mem_reg_156__7_ ( .D(n5855), .CK(clk), .Q(n[1360]), .QN(n1937) );
  DFF_X1 reg_mem_reg_156__6_ ( .D(n5854), .CK(clk), .Q(n[1359]), .QN(n1938) );
  DFF_X1 reg_mem_reg_156__5_ ( .D(n5853), .CK(clk), .Q(n[1358]), .QN(n1939) );
  DFF_X1 reg_mem_reg_156__4_ ( .D(n5852), .CK(clk), .Q(n[1357]), .QN(n1940) );
  DFF_X1 reg_mem_reg_156__3_ ( .D(n5851), .CK(clk), .Q(n[1356]), .QN(n1941) );
  DFF_X1 reg_mem_reg_156__2_ ( .D(n5850), .CK(clk), .Q(n[1355]), .QN(n1942) );
  DFF_X1 reg_mem_reg_156__1_ ( .D(n5849), .CK(clk), .Q(n[1354]), .QN(n1943) );
  DFF_X1 reg_mem_reg_156__0_ ( .D(n5848), .CK(clk), .Q(n[1353]), .QN(n1944) );
  DFF_X1 reg_mem_reg_157__7_ ( .D(n5847), .CK(clk), .Q(n[1352]), .QN(n1945) );
  DFF_X1 reg_mem_reg_157__6_ ( .D(n5846), .CK(clk), .Q(n[1351]), .QN(n1946) );
  DFF_X1 reg_mem_reg_157__5_ ( .D(n5845), .CK(clk), .Q(n[1350]), .QN(n1947) );
  DFF_X1 reg_mem_reg_157__4_ ( .D(n5844), .CK(clk), .Q(n[1349]), .QN(n1948) );
  DFF_X1 reg_mem_reg_157__3_ ( .D(n5843), .CK(clk), .Q(n[1348]), .QN(n1949) );
  DFF_X1 reg_mem_reg_157__2_ ( .D(n5842), .CK(clk), .Q(n[1347]), .QN(n1950) );
  DFF_X1 reg_mem_reg_157__1_ ( .D(n5841), .CK(clk), .Q(n[1346]), .QN(n1951) );
  DFF_X1 reg_mem_reg_157__0_ ( .D(n5840), .CK(clk), .Q(n[1345]), .QN(n1952) );
  DFF_X1 reg_mem_reg_158__7_ ( .D(n5839), .CK(clk), .QN(n1969) );
  DFF_X1 reg_mem_reg_158__6_ ( .D(n5838), .CK(clk), .QN(n1970) );
  DFF_X1 reg_mem_reg_158__5_ ( .D(n5837), .CK(clk), .QN(n1971) );
  DFF_X1 reg_mem_reg_158__4_ ( .D(n5836), .CK(clk), .QN(n1972) );
  DFF_X1 reg_mem_reg_158__3_ ( .D(n5835), .CK(clk), .QN(n1973) );
  DFF_X1 reg_mem_reg_158__2_ ( .D(n5834), .CK(clk), .QN(n1974) );
  DFF_X1 reg_mem_reg_158__1_ ( .D(n5833), .CK(clk), .QN(n1975) );
  DFF_X1 reg_mem_reg_158__0_ ( .D(n5832), .CK(clk), .QN(n1976) );
  DFF_X1 reg_mem_reg_159__7_ ( .D(n5831), .CK(clk), .QN(n1977) );
  DFF_X1 reg_mem_reg_159__6_ ( .D(n5830), .CK(clk), .QN(n1978) );
  DFF_X1 reg_mem_reg_159__5_ ( .D(n5829), .CK(clk), .QN(n1979) );
  DFF_X1 reg_mem_reg_159__4_ ( .D(n5828), .CK(clk), .QN(n1980) );
  DFF_X1 reg_mem_reg_159__3_ ( .D(n5827), .CK(clk), .QN(n1981) );
  DFF_X1 reg_mem_reg_159__2_ ( .D(n5826), .CK(clk), .QN(n1982) );
  DFF_X1 reg_mem_reg_159__1_ ( .D(n5825), .CK(clk), .QN(n1983) );
  DFF_X1 reg_mem_reg_159__0_ ( .D(n5824), .CK(clk), .QN(n1984) );
  DFF_X1 reg_mem_reg_160__7_ ( .D(n5823), .CK(clk), .Q(n[1328]), .QN(n2001) );
  DFF_X1 reg_mem_reg_160__6_ ( .D(n5822), .CK(clk), .Q(n[1327]), .QN(n2002) );
  DFF_X1 reg_mem_reg_160__5_ ( .D(n5821), .CK(clk), .Q(n[1326]), .QN(n2003) );
  DFF_X1 reg_mem_reg_160__4_ ( .D(n5820), .CK(clk), .Q(n[1325]), .QN(n2004) );
  DFF_X1 reg_mem_reg_160__3_ ( .D(n5819), .CK(clk), .Q(n[1324]), .QN(n2005) );
  DFF_X1 reg_mem_reg_160__2_ ( .D(n5818), .CK(clk), .Q(n[1323]), .QN(n2006) );
  DFF_X1 reg_mem_reg_160__1_ ( .D(n5817), .CK(clk), .Q(n[1322]), .QN(n2007) );
  DFF_X1 reg_mem_reg_160__0_ ( .D(n5816), .CK(clk), .Q(n[1321]), .QN(n2008) );
  DFF_X1 reg_mem_reg_161__7_ ( .D(n5815), .CK(clk), .Q(n[1320]), .QN(n2009) );
  DFF_X1 reg_mem_reg_161__6_ ( .D(n5814), .CK(clk), .Q(n[1319]), .QN(n2010) );
  DFF_X1 reg_mem_reg_161__5_ ( .D(n5813), .CK(clk), .Q(n[1318]), .QN(n2011) );
  DFF_X1 reg_mem_reg_161__4_ ( .D(n5812), .CK(clk), .Q(n[1317]), .QN(n2012) );
  DFF_X1 reg_mem_reg_161__3_ ( .D(n5811), .CK(clk), .Q(n[1316]), .QN(n2013) );
  DFF_X1 reg_mem_reg_161__2_ ( .D(n5810), .CK(clk), .Q(n[1315]), .QN(n2014) );
  DFF_X1 reg_mem_reg_161__1_ ( .D(n5809), .CK(clk), .Q(n[1314]), .QN(n2015) );
  DFF_X1 reg_mem_reg_161__0_ ( .D(n5808), .CK(clk), .Q(n[1313]), .QN(n2016) );
  DFF_X1 reg_mem_reg_162__7_ ( .D(n5807), .CK(clk), .QN(n2033) );
  DFF_X1 reg_mem_reg_162__6_ ( .D(n5806), .CK(clk), .QN(n2034) );
  DFF_X1 reg_mem_reg_162__5_ ( .D(n5805), .CK(clk), .QN(n2035) );
  DFF_X1 reg_mem_reg_162__4_ ( .D(n5804), .CK(clk), .QN(n2036) );
  DFF_X1 reg_mem_reg_162__3_ ( .D(n5803), .CK(clk), .QN(n2037) );
  DFF_X1 reg_mem_reg_162__2_ ( .D(n5802), .CK(clk), .QN(n2038) );
  DFF_X1 reg_mem_reg_162__1_ ( .D(n5801), .CK(clk), .QN(n2039) );
  DFF_X1 reg_mem_reg_162__0_ ( .D(n5800), .CK(clk), .QN(n2040) );
  DFF_X1 reg_mem_reg_163__7_ ( .D(n5799), .CK(clk), .QN(n2041) );
  DFF_X1 reg_mem_reg_163__6_ ( .D(n5798), .CK(clk), .QN(n2042) );
  DFF_X1 reg_mem_reg_163__5_ ( .D(n5797), .CK(clk), .QN(n2043) );
  DFF_X1 reg_mem_reg_163__4_ ( .D(n5796), .CK(clk), .QN(n2044) );
  DFF_X1 reg_mem_reg_163__3_ ( .D(n5795), .CK(clk), .QN(n2045) );
  DFF_X1 reg_mem_reg_163__2_ ( .D(n5794), .CK(clk), .QN(n2046) );
  DFF_X1 reg_mem_reg_163__1_ ( .D(n5793), .CK(clk), .QN(n2047) );
  DFF_X1 reg_mem_reg_163__0_ ( .D(n5792), .CK(clk), .QN(n2048) );
  DFF_X1 reg_mem_reg_164__7_ ( .D(n5791), .CK(clk), .Q(n[1296]), .QN(n2065) );
  DFF_X1 reg_mem_reg_164__6_ ( .D(n5790), .CK(clk), .Q(n[1295]), .QN(n2066) );
  DFF_X1 reg_mem_reg_164__5_ ( .D(n5789), .CK(clk), .Q(n[1294]), .QN(n2067) );
  DFF_X1 reg_mem_reg_164__4_ ( .D(n5788), .CK(clk), .Q(n[1293]), .QN(n2068) );
  DFF_X1 reg_mem_reg_164__3_ ( .D(n5787), .CK(clk), .Q(n[1292]), .QN(n2069) );
  DFF_X1 reg_mem_reg_164__2_ ( .D(n5786), .CK(clk), .Q(n[1291]), .QN(n2070) );
  DFF_X1 reg_mem_reg_164__1_ ( .D(n5785), .CK(clk), .Q(n[1290]), .QN(n2071) );
  DFF_X1 reg_mem_reg_164__0_ ( .D(n5784), .CK(clk), .Q(n[1289]), .QN(n2072) );
  DFF_X1 reg_mem_reg_165__7_ ( .D(n5783), .CK(clk), .Q(n[1288]), .QN(n2073) );
  DFF_X1 reg_mem_reg_165__6_ ( .D(n5782), .CK(clk), .Q(n[1287]), .QN(n2074) );
  DFF_X1 reg_mem_reg_165__5_ ( .D(n5781), .CK(clk), .Q(n[1286]), .QN(n2075) );
  DFF_X1 reg_mem_reg_165__4_ ( .D(n5780), .CK(clk), .Q(n[1285]), .QN(n2076) );
  DFF_X1 reg_mem_reg_165__3_ ( .D(n5779), .CK(clk), .Q(n[1284]), .QN(n2077) );
  DFF_X1 reg_mem_reg_165__2_ ( .D(n5778), .CK(clk), .Q(n[1283]), .QN(n2078) );
  DFF_X1 reg_mem_reg_165__1_ ( .D(n5777), .CK(clk), .Q(n[1282]), .QN(n2079) );
  DFF_X1 reg_mem_reg_165__0_ ( .D(n5776), .CK(clk), .Q(n[1281]), .QN(n2080) );
  DFF_X1 reg_mem_reg_166__7_ ( .D(n5775), .CK(clk), .QN(n2097) );
  DFF_X1 reg_mem_reg_166__6_ ( .D(n5774), .CK(clk), .QN(n2098) );
  DFF_X1 reg_mem_reg_166__5_ ( .D(n5773), .CK(clk), .QN(n2099) );
  DFF_X1 reg_mem_reg_166__4_ ( .D(n5772), .CK(clk), .QN(n2100) );
  DFF_X1 reg_mem_reg_166__3_ ( .D(n5771), .CK(clk), .QN(n2101) );
  DFF_X1 reg_mem_reg_166__2_ ( .D(n5770), .CK(clk), .QN(n2102) );
  DFF_X1 reg_mem_reg_166__1_ ( .D(n5769), .CK(clk), .QN(n2103) );
  DFF_X1 reg_mem_reg_166__0_ ( .D(n5768), .CK(clk), .QN(n2104) );
  DFF_X1 reg_mem_reg_167__7_ ( .D(n5767), .CK(clk), .QN(n2105) );
  DFF_X1 reg_mem_reg_167__6_ ( .D(n5766), .CK(clk), .QN(n2106) );
  DFF_X1 reg_mem_reg_167__5_ ( .D(n5765), .CK(clk), .QN(n2107) );
  DFF_X1 reg_mem_reg_167__4_ ( .D(n5764), .CK(clk), .QN(n2108) );
  DFF_X1 reg_mem_reg_167__3_ ( .D(n5763), .CK(clk), .QN(n2109) );
  DFF_X1 reg_mem_reg_167__2_ ( .D(n5762), .CK(clk), .QN(n2110) );
  DFF_X1 reg_mem_reg_167__1_ ( .D(n5761), .CK(clk), .QN(n2111) );
  DFF_X1 reg_mem_reg_167__0_ ( .D(n5760), .CK(clk), .QN(n2112) );
  DFF_X1 reg_mem_reg_168__7_ ( .D(n5759), .CK(clk), .Q(n[1264]), .QN(n2129) );
  DFF_X1 reg_mem_reg_168__6_ ( .D(n5758), .CK(clk), .Q(n[1263]), .QN(n2130) );
  DFF_X1 reg_mem_reg_168__5_ ( .D(n5757), .CK(clk), .Q(n[1262]), .QN(n2131) );
  DFF_X1 reg_mem_reg_168__4_ ( .D(n5756), .CK(clk), .Q(n[1261]), .QN(n2132) );
  DFF_X1 reg_mem_reg_168__3_ ( .D(n5755), .CK(clk), .Q(n[1260]), .QN(n2133) );
  DFF_X1 reg_mem_reg_168__2_ ( .D(n5754), .CK(clk), .Q(n[1259]), .QN(n2134) );
  DFF_X1 reg_mem_reg_168__1_ ( .D(n5753), .CK(clk), .Q(n[1258]), .QN(n2135) );
  DFF_X1 reg_mem_reg_168__0_ ( .D(n5752), .CK(clk), .Q(n[1257]), .QN(n2136) );
  DFF_X1 reg_mem_reg_169__7_ ( .D(n5751), .CK(clk), .Q(n[1256]), .QN(n2137) );
  DFF_X1 reg_mem_reg_169__6_ ( .D(n5750), .CK(clk), .Q(n[1255]), .QN(n2138) );
  DFF_X1 reg_mem_reg_169__5_ ( .D(n5749), .CK(clk), .Q(n[1254]), .QN(n2139) );
  DFF_X1 reg_mem_reg_169__4_ ( .D(n5748), .CK(clk), .Q(n[1253]), .QN(n2140) );
  DFF_X1 reg_mem_reg_169__3_ ( .D(n5747), .CK(clk), .Q(n[1252]), .QN(n2141) );
  DFF_X1 reg_mem_reg_169__2_ ( .D(n5746), .CK(clk), .Q(n[1251]), .QN(n2142) );
  DFF_X1 reg_mem_reg_169__1_ ( .D(n5745), .CK(clk), .Q(n[1250]), .QN(n2143) );
  DFF_X1 reg_mem_reg_169__0_ ( .D(n5744), .CK(clk), .Q(n[1249]), .QN(n2144) );
  DFF_X1 reg_mem_reg_170__7_ ( .D(n5743), .CK(clk), .QN(n2161) );
  DFF_X1 reg_mem_reg_170__6_ ( .D(n5742), .CK(clk), .QN(n2162) );
  DFF_X1 reg_mem_reg_170__5_ ( .D(n5741), .CK(clk), .QN(n2163) );
  DFF_X1 reg_mem_reg_170__4_ ( .D(n5740), .CK(clk), .QN(n2164) );
  DFF_X1 reg_mem_reg_170__3_ ( .D(n5739), .CK(clk), .QN(n2165) );
  DFF_X1 reg_mem_reg_170__2_ ( .D(n5738), .CK(clk), .QN(n2166) );
  DFF_X1 reg_mem_reg_170__1_ ( .D(n5737), .CK(clk), .QN(n2167) );
  DFF_X1 reg_mem_reg_170__0_ ( .D(n5736), .CK(clk), .QN(n2168) );
  DFF_X1 reg_mem_reg_171__7_ ( .D(n5735), .CK(clk), .QN(n2169) );
  DFF_X1 reg_mem_reg_171__6_ ( .D(n5734), .CK(clk), .QN(n2170) );
  DFF_X1 reg_mem_reg_171__5_ ( .D(n5733), .CK(clk), .QN(n2171) );
  DFF_X1 reg_mem_reg_171__4_ ( .D(n5732), .CK(clk), .QN(n2172) );
  DFF_X1 reg_mem_reg_171__3_ ( .D(n5731), .CK(clk), .QN(n2173) );
  DFF_X1 reg_mem_reg_171__2_ ( .D(n5730), .CK(clk), .QN(n2174) );
  DFF_X1 reg_mem_reg_171__1_ ( .D(n5729), .CK(clk), .QN(n2175) );
  DFF_X1 reg_mem_reg_171__0_ ( .D(n5728), .CK(clk), .QN(n2176) );
  DFF_X1 reg_mem_reg_172__7_ ( .D(n5727), .CK(clk), .Q(n[1232]), .QN(n2193) );
  DFF_X1 reg_mem_reg_172__6_ ( .D(n5726), .CK(clk), .Q(n[1231]), .QN(n2194) );
  DFF_X1 reg_mem_reg_172__5_ ( .D(n5725), .CK(clk), .Q(n[1230]), .QN(n2195) );
  DFF_X1 reg_mem_reg_172__4_ ( .D(n5724), .CK(clk), .Q(n[1229]), .QN(n2196) );
  DFF_X1 reg_mem_reg_172__3_ ( .D(n5723), .CK(clk), .Q(n[1228]), .QN(n2197) );
  DFF_X1 reg_mem_reg_172__2_ ( .D(n5722), .CK(clk), .Q(n[1227]), .QN(n2198) );
  DFF_X1 reg_mem_reg_172__1_ ( .D(n5721), .CK(clk), .Q(n[1226]), .QN(n2199) );
  DFF_X1 reg_mem_reg_172__0_ ( .D(n5720), .CK(clk), .Q(n[1225]), .QN(n2200) );
  DFF_X1 reg_mem_reg_173__7_ ( .D(n5719), .CK(clk), .Q(n[1224]), .QN(n2201) );
  DFF_X1 reg_mem_reg_173__6_ ( .D(n5718), .CK(clk), .Q(n[1223]), .QN(n2202) );
  DFF_X1 reg_mem_reg_173__5_ ( .D(n5717), .CK(clk), .Q(n[1222]), .QN(n2203) );
  DFF_X1 reg_mem_reg_173__4_ ( .D(n5716), .CK(clk), .Q(n[1221]), .QN(n2204) );
  DFF_X1 reg_mem_reg_173__3_ ( .D(n5715), .CK(clk), .Q(n[1220]), .QN(n2205) );
  DFF_X1 reg_mem_reg_173__2_ ( .D(n5714), .CK(clk), .Q(n[1219]), .QN(n2206) );
  DFF_X1 reg_mem_reg_173__1_ ( .D(n5713), .CK(clk), .Q(n[1218]), .QN(n2207) );
  DFF_X1 reg_mem_reg_173__0_ ( .D(n5712), .CK(clk), .Q(n[1217]), .QN(n2208) );
  DFF_X1 reg_mem_reg_174__7_ ( .D(n5711), .CK(clk), .QN(n2225) );
  DFF_X1 reg_mem_reg_174__6_ ( .D(n5710), .CK(clk), .QN(n2226) );
  DFF_X1 reg_mem_reg_174__5_ ( .D(n5709), .CK(clk), .QN(n2227) );
  DFF_X1 reg_mem_reg_174__4_ ( .D(n5708), .CK(clk), .QN(n2228) );
  DFF_X1 reg_mem_reg_174__3_ ( .D(n5707), .CK(clk), .QN(n2229) );
  DFF_X1 reg_mem_reg_174__2_ ( .D(n5706), .CK(clk), .QN(n2230) );
  DFF_X1 reg_mem_reg_174__1_ ( .D(n5705), .CK(clk), .QN(n2231) );
  DFF_X1 reg_mem_reg_174__0_ ( .D(n5704), .CK(clk), .QN(n2232) );
  DFF_X1 reg_mem_reg_175__7_ ( .D(n5703), .CK(clk), .QN(n2233) );
  DFF_X1 reg_mem_reg_175__6_ ( .D(n5702), .CK(clk), .QN(n2234) );
  DFF_X1 reg_mem_reg_175__5_ ( .D(n5701), .CK(clk), .QN(n2235) );
  DFF_X1 reg_mem_reg_175__4_ ( .D(n5700), .CK(clk), .QN(n2236) );
  DFF_X1 reg_mem_reg_175__3_ ( .D(n5699), .CK(clk), .QN(n2237) );
  DFF_X1 reg_mem_reg_175__2_ ( .D(n5698), .CK(clk), .QN(n2238) );
  DFF_X1 reg_mem_reg_175__1_ ( .D(n5697), .CK(clk), .QN(n2239) );
  DFF_X1 reg_mem_reg_175__0_ ( .D(n5696), .CK(clk), .QN(n2240) );
  DFF_X1 reg_mem_reg_176__7_ ( .D(n5695), .CK(clk), .Q(n[1200]), .QN(n2257) );
  DFF_X1 reg_mem_reg_176__6_ ( .D(n5694), .CK(clk), .Q(n[1199]), .QN(n2258) );
  DFF_X1 reg_mem_reg_176__5_ ( .D(n5693), .CK(clk), .Q(n[1198]), .QN(n2259) );
  DFF_X1 reg_mem_reg_176__4_ ( .D(n5692), .CK(clk), .Q(n[1197]), .QN(n2260) );
  DFF_X1 reg_mem_reg_176__3_ ( .D(n5691), .CK(clk), .Q(n[1196]), .QN(n2261) );
  DFF_X1 reg_mem_reg_176__2_ ( .D(n5690), .CK(clk), .Q(n[1195]), .QN(n2262) );
  DFF_X1 reg_mem_reg_176__1_ ( .D(n5689), .CK(clk), .Q(n[1194]), .QN(n2263) );
  DFF_X1 reg_mem_reg_176__0_ ( .D(n5688), .CK(clk), .Q(n[1193]), .QN(n2264) );
  DFF_X1 reg_mem_reg_177__7_ ( .D(n5687), .CK(clk), .Q(n[1192]), .QN(n2265) );
  DFF_X1 reg_mem_reg_177__6_ ( .D(n5686), .CK(clk), .Q(n[1191]), .QN(n2266) );
  DFF_X1 reg_mem_reg_177__5_ ( .D(n5685), .CK(clk), .Q(n[1190]), .QN(n2267) );
  DFF_X1 reg_mem_reg_177__4_ ( .D(n5684), .CK(clk), .Q(n[1189]), .QN(n2268) );
  DFF_X1 reg_mem_reg_177__3_ ( .D(n5683), .CK(clk), .Q(n[1188]), .QN(n2269) );
  DFF_X1 reg_mem_reg_177__2_ ( .D(n5682), .CK(clk), .Q(n[1187]), .QN(n2270) );
  DFF_X1 reg_mem_reg_177__1_ ( .D(n5681), .CK(clk), .Q(n[1186]), .QN(n2271) );
  DFF_X1 reg_mem_reg_177__0_ ( .D(n5680), .CK(clk), .Q(n[1185]), .QN(n2272) );
  DFF_X1 reg_mem_reg_178__7_ ( .D(n5679), .CK(clk), .QN(n2289) );
  DFF_X1 reg_mem_reg_178__6_ ( .D(n5678), .CK(clk), .QN(n2290) );
  DFF_X1 reg_mem_reg_178__5_ ( .D(n5677), .CK(clk), .QN(n2291) );
  DFF_X1 reg_mem_reg_178__4_ ( .D(n5676), .CK(clk), .QN(n2292) );
  DFF_X1 reg_mem_reg_178__3_ ( .D(n5675), .CK(clk), .QN(n2293) );
  DFF_X1 reg_mem_reg_178__2_ ( .D(n5674), .CK(clk), .QN(n2294) );
  DFF_X1 reg_mem_reg_178__1_ ( .D(n5673), .CK(clk), .QN(n2295) );
  DFF_X1 reg_mem_reg_178__0_ ( .D(n5672), .CK(clk), .QN(n2296) );
  DFF_X1 reg_mem_reg_179__7_ ( .D(n5671), .CK(clk), .QN(n2297) );
  DFF_X1 reg_mem_reg_179__6_ ( .D(n5670), .CK(clk), .QN(n2298) );
  DFF_X1 reg_mem_reg_179__5_ ( .D(n5669), .CK(clk), .QN(n2299) );
  DFF_X1 reg_mem_reg_179__4_ ( .D(n5668), .CK(clk), .QN(n2300) );
  DFF_X1 reg_mem_reg_179__3_ ( .D(n5667), .CK(clk), .QN(n2301) );
  DFF_X1 reg_mem_reg_179__2_ ( .D(n5666), .CK(clk), .QN(n2302) );
  DFF_X1 reg_mem_reg_179__1_ ( .D(n5665), .CK(clk), .QN(n2303) );
  DFF_X1 reg_mem_reg_179__0_ ( .D(n5664), .CK(clk), .QN(n2304) );
  DFF_X1 reg_mem_reg_180__7_ ( .D(n5663), .CK(clk), .Q(n[1168]), .QN(n2321) );
  DFF_X1 reg_mem_reg_180__6_ ( .D(n5662), .CK(clk), .Q(n[1167]), .QN(n2322) );
  DFF_X1 reg_mem_reg_180__5_ ( .D(n5661), .CK(clk), .Q(n[1166]), .QN(n2323) );
  DFF_X1 reg_mem_reg_180__4_ ( .D(n5660), .CK(clk), .Q(n[1165]), .QN(n2324) );
  DFF_X1 reg_mem_reg_180__3_ ( .D(n5659), .CK(clk), .Q(n[1164]), .QN(n2325) );
  DFF_X1 reg_mem_reg_180__2_ ( .D(n5658), .CK(clk), .Q(n[1163]), .QN(n2326) );
  DFF_X1 reg_mem_reg_180__1_ ( .D(n5657), .CK(clk), .Q(n[1162]), .QN(n2327) );
  DFF_X1 reg_mem_reg_180__0_ ( .D(n5656), .CK(clk), .Q(n[1161]), .QN(n2328) );
  DFF_X1 reg_mem_reg_181__7_ ( .D(n5655), .CK(clk), .Q(n[1160]), .QN(n2329) );
  DFF_X1 reg_mem_reg_181__6_ ( .D(n5654), .CK(clk), .Q(n[1159]), .QN(n2330) );
  DFF_X1 reg_mem_reg_181__5_ ( .D(n5653), .CK(clk), .Q(n[1158]), .QN(n2331) );
  DFF_X1 reg_mem_reg_181__4_ ( .D(n5652), .CK(clk), .Q(n[1157]), .QN(n2332) );
  DFF_X1 reg_mem_reg_181__3_ ( .D(n5651), .CK(clk), .Q(n[1156]), .QN(n2333) );
  DFF_X1 reg_mem_reg_181__2_ ( .D(n5650), .CK(clk), .Q(n[1155]), .QN(n2334) );
  DFF_X1 reg_mem_reg_181__1_ ( .D(n5649), .CK(clk), .Q(n[1154]), .QN(n2335) );
  DFF_X1 reg_mem_reg_181__0_ ( .D(n5648), .CK(clk), .Q(n[1153]), .QN(n2336) );
  DFF_X1 reg_mem_reg_182__7_ ( .D(n5647), .CK(clk), .QN(n2353) );
  DFF_X1 reg_mem_reg_182__6_ ( .D(n5646), .CK(clk), .QN(n2354) );
  DFF_X1 reg_mem_reg_182__5_ ( .D(n5645), .CK(clk), .QN(n2355) );
  DFF_X1 reg_mem_reg_182__4_ ( .D(n5644), .CK(clk), .QN(n2356) );
  DFF_X1 reg_mem_reg_182__3_ ( .D(n5643), .CK(clk), .QN(n2357) );
  DFF_X1 reg_mem_reg_182__2_ ( .D(n5642), .CK(clk), .QN(n2358) );
  DFF_X1 reg_mem_reg_182__1_ ( .D(n5641), .CK(clk), .QN(n2359) );
  DFF_X1 reg_mem_reg_182__0_ ( .D(n5640), .CK(clk), .QN(n2360) );
  DFF_X1 reg_mem_reg_183__7_ ( .D(n5639), .CK(clk), .QN(n2361) );
  DFF_X1 reg_mem_reg_183__6_ ( .D(n5638), .CK(clk), .QN(n2362) );
  DFF_X1 reg_mem_reg_183__5_ ( .D(n5637), .CK(clk), .QN(n2363) );
  DFF_X1 reg_mem_reg_183__4_ ( .D(n5636), .CK(clk), .QN(n2364) );
  DFF_X1 reg_mem_reg_183__3_ ( .D(n5635), .CK(clk), .QN(n2365) );
  DFF_X1 reg_mem_reg_183__2_ ( .D(n5634), .CK(clk), .QN(n2366) );
  DFF_X1 reg_mem_reg_183__1_ ( .D(n5633), .CK(clk), .QN(n2367) );
  DFF_X1 reg_mem_reg_183__0_ ( .D(n5632), .CK(clk), .QN(n2368) );
  DFF_X1 reg_mem_reg_184__7_ ( .D(n5631), .CK(clk), .Q(n[1136]), .QN(n2385) );
  DFF_X1 reg_mem_reg_184__6_ ( .D(n5630), .CK(clk), .Q(n[1135]), .QN(n2386) );
  DFF_X1 reg_mem_reg_184__5_ ( .D(n5629), .CK(clk), .Q(n[1134]), .QN(n2387) );
  DFF_X1 reg_mem_reg_184__4_ ( .D(n5628), .CK(clk), .Q(n[1133]), .QN(n2388) );
  DFF_X1 reg_mem_reg_184__3_ ( .D(n5627), .CK(clk), .Q(n[1132]), .QN(n2389) );
  DFF_X1 reg_mem_reg_184__2_ ( .D(n5626), .CK(clk), .Q(n[1131]), .QN(n2390) );
  DFF_X1 reg_mem_reg_184__1_ ( .D(n5625), .CK(clk), .Q(n[1130]), .QN(n2391) );
  DFF_X1 reg_mem_reg_184__0_ ( .D(n5624), .CK(clk), .Q(n[1129]), .QN(n2392) );
  DFF_X1 reg_mem_reg_185__7_ ( .D(n5623), .CK(clk), .Q(n[1128]), .QN(n2393) );
  DFF_X1 reg_mem_reg_185__6_ ( .D(n5622), .CK(clk), .Q(n[1127]), .QN(n2394) );
  DFF_X1 reg_mem_reg_185__5_ ( .D(n5621), .CK(clk), .Q(n[1126]), .QN(n2395) );
  DFF_X1 reg_mem_reg_185__4_ ( .D(n5620), .CK(clk), .Q(n[1125]), .QN(n2396) );
  DFF_X1 reg_mem_reg_185__3_ ( .D(n5619), .CK(clk), .Q(n[1124]), .QN(n2397) );
  DFF_X1 reg_mem_reg_185__2_ ( .D(n5618), .CK(clk), .Q(n[1123]), .QN(n2398) );
  DFF_X1 reg_mem_reg_185__1_ ( .D(n5617), .CK(clk), .Q(n[1122]), .QN(n2399) );
  DFF_X1 reg_mem_reg_185__0_ ( .D(n5616), .CK(clk), .Q(n[1121]), .QN(n2400) );
  DFF_X1 reg_mem_reg_186__7_ ( .D(n5615), .CK(clk), .QN(n2417) );
  DFF_X1 reg_mem_reg_186__6_ ( .D(n5614), .CK(clk), .QN(n2418) );
  DFF_X1 reg_mem_reg_186__5_ ( .D(n5613), .CK(clk), .QN(n2419) );
  DFF_X1 reg_mem_reg_186__4_ ( .D(n5612), .CK(clk), .QN(n2420) );
  DFF_X1 reg_mem_reg_186__3_ ( .D(n5611), .CK(clk), .QN(n2421) );
  DFF_X1 reg_mem_reg_186__2_ ( .D(n5610), .CK(clk), .QN(n2422) );
  DFF_X1 reg_mem_reg_186__1_ ( .D(n5609), .CK(clk), .QN(n2423) );
  DFF_X1 reg_mem_reg_186__0_ ( .D(n5608), .CK(clk), .QN(n2424) );
  DFF_X1 reg_mem_reg_187__7_ ( .D(n5607), .CK(clk), .QN(n2425) );
  DFF_X1 reg_mem_reg_187__6_ ( .D(n5606), .CK(clk), .QN(n2426) );
  DFF_X1 reg_mem_reg_187__5_ ( .D(n5605), .CK(clk), .QN(n2427) );
  DFF_X1 reg_mem_reg_187__4_ ( .D(n5604), .CK(clk), .QN(n2428) );
  DFF_X1 reg_mem_reg_187__3_ ( .D(n5603), .CK(clk), .QN(n2429) );
  DFF_X1 reg_mem_reg_187__2_ ( .D(n5602), .CK(clk), .QN(n2430) );
  DFF_X1 reg_mem_reg_187__1_ ( .D(n5601), .CK(clk), .QN(n2431) );
  DFF_X1 reg_mem_reg_187__0_ ( .D(n5600), .CK(clk), .QN(n2432) );
  DFF_X1 reg_mem_reg_188__7_ ( .D(n5599), .CK(clk), .Q(n[1104]), .QN(n2449) );
  DFF_X1 reg_mem_reg_188__6_ ( .D(n5598), .CK(clk), .Q(n[1103]), .QN(n2450) );
  DFF_X1 reg_mem_reg_188__5_ ( .D(n5597), .CK(clk), .Q(n[1102]), .QN(n2451) );
  DFF_X1 reg_mem_reg_188__4_ ( .D(n5596), .CK(clk), .Q(n[1101]), .QN(n2452) );
  DFF_X1 reg_mem_reg_188__3_ ( .D(n5595), .CK(clk), .Q(n[1100]), .QN(n2453) );
  DFF_X1 reg_mem_reg_188__2_ ( .D(n5594), .CK(clk), .Q(n[1099]), .QN(n2454) );
  DFF_X1 reg_mem_reg_188__1_ ( .D(n5593), .CK(clk), .Q(n[1098]), .QN(n2455) );
  DFF_X1 reg_mem_reg_188__0_ ( .D(n5592), .CK(clk), .Q(n[1097]), .QN(n2456) );
  DFF_X1 reg_mem_reg_189__7_ ( .D(n5591), .CK(clk), .Q(n[1096]), .QN(n2457) );
  DFF_X1 reg_mem_reg_189__6_ ( .D(n5590), .CK(clk), .Q(n[1095]), .QN(n2458) );
  DFF_X1 reg_mem_reg_189__5_ ( .D(n5589), .CK(clk), .Q(n[1094]), .QN(n2459) );
  DFF_X1 reg_mem_reg_189__4_ ( .D(n5588), .CK(clk), .Q(n[1093]), .QN(n2460) );
  DFF_X1 reg_mem_reg_189__3_ ( .D(n5587), .CK(clk), .Q(n[1092]), .QN(n2461) );
  DFF_X1 reg_mem_reg_189__2_ ( .D(n5586), .CK(clk), .Q(n[1091]), .QN(n2462) );
  DFF_X1 reg_mem_reg_189__1_ ( .D(n5585), .CK(clk), .Q(n[1090]), .QN(n2463) );
  DFF_X1 reg_mem_reg_189__0_ ( .D(n5584), .CK(clk), .Q(n[1089]), .QN(n2464) );
  DFF_X1 reg_mem_reg_190__7_ ( .D(n5583), .CK(clk), .QN(n2481) );
  DFF_X1 reg_mem_reg_190__6_ ( .D(n5582), .CK(clk), .QN(n2482) );
  DFF_X1 reg_mem_reg_190__5_ ( .D(n5581), .CK(clk), .QN(n2483) );
  DFF_X1 reg_mem_reg_190__4_ ( .D(n5580), .CK(clk), .QN(n2484) );
  DFF_X1 reg_mem_reg_190__3_ ( .D(n5579), .CK(clk), .QN(n2485) );
  DFF_X1 reg_mem_reg_190__2_ ( .D(n5578), .CK(clk), .QN(n2486) );
  DFF_X1 reg_mem_reg_190__1_ ( .D(n5577), .CK(clk), .QN(n2487) );
  DFF_X1 reg_mem_reg_190__0_ ( .D(n5576), .CK(clk), .QN(n2488) );
  DFF_X1 reg_mem_reg_191__7_ ( .D(n5575), .CK(clk), .QN(n2489) );
  DFF_X1 reg_mem_reg_191__6_ ( .D(n5574), .CK(clk), .QN(n2490) );
  DFF_X1 reg_mem_reg_191__5_ ( .D(n5573), .CK(clk), .QN(n2491) );
  DFF_X1 reg_mem_reg_191__4_ ( .D(n5572), .CK(clk), .QN(n2492) );
  DFF_X1 reg_mem_reg_191__3_ ( .D(n5571), .CK(clk), .QN(n2493) );
  DFF_X1 reg_mem_reg_191__2_ ( .D(n5570), .CK(clk), .QN(n2494) );
  DFF_X1 reg_mem_reg_191__1_ ( .D(n5569), .CK(clk), .QN(n2495) );
  DFF_X1 reg_mem_reg_191__0_ ( .D(n5568), .CK(clk), .QN(n2496) );
  DFF_X1 reg_mem_reg_192__7_ ( .D(n5567), .CK(clk), .Q(n[1072]), .QN(n2513) );
  DFF_X1 reg_mem_reg_192__6_ ( .D(n5566), .CK(clk), .Q(n[1071]), .QN(n2514) );
  DFF_X1 reg_mem_reg_192__5_ ( .D(n5565), .CK(clk), .Q(n[1070]), .QN(n2515) );
  DFF_X1 reg_mem_reg_192__4_ ( .D(n5564), .CK(clk), .Q(n[1069]), .QN(n2516) );
  DFF_X1 reg_mem_reg_192__3_ ( .D(n5563), .CK(clk), .Q(n[1068]), .QN(n2517) );
  DFF_X1 reg_mem_reg_192__2_ ( .D(n5562), .CK(clk), .Q(n[1067]), .QN(n2518) );
  DFF_X1 reg_mem_reg_192__1_ ( .D(n5561), .CK(clk), .Q(n[1066]), .QN(n2519) );
  DFF_X1 reg_mem_reg_192__0_ ( .D(n5560), .CK(clk), .Q(n[1065]), .QN(n2520) );
  DFF_X1 reg_mem_reg_193__7_ ( .D(n5559), .CK(clk), .Q(n[1064]), .QN(n2521) );
  DFF_X1 reg_mem_reg_193__6_ ( .D(n5558), .CK(clk), .Q(n[1063]), .QN(n2522) );
  DFF_X1 reg_mem_reg_193__5_ ( .D(n5557), .CK(clk), .Q(n[1062]), .QN(n2523) );
  DFF_X1 reg_mem_reg_193__4_ ( .D(n5556), .CK(clk), .Q(n[1061]), .QN(n2524) );
  DFF_X1 reg_mem_reg_193__3_ ( .D(n5555), .CK(clk), .Q(n[1060]), .QN(n2525) );
  DFF_X1 reg_mem_reg_193__2_ ( .D(n5554), .CK(clk), .Q(n[1059]), .QN(n2526) );
  DFF_X1 reg_mem_reg_193__1_ ( .D(n5553), .CK(clk), .Q(n[1058]), .QN(n2527) );
  DFF_X1 reg_mem_reg_193__0_ ( .D(n5552), .CK(clk), .Q(n[1057]), .QN(n2528) );
  DFF_X1 reg_mem_reg_194__7_ ( .D(n5551), .CK(clk), .QN(n2545) );
  DFF_X1 reg_mem_reg_194__6_ ( .D(n5550), .CK(clk), .QN(n2546) );
  DFF_X1 reg_mem_reg_194__5_ ( .D(n5549), .CK(clk), .QN(n2547) );
  DFF_X1 reg_mem_reg_194__4_ ( .D(n5548), .CK(clk), .QN(n2548) );
  DFF_X1 reg_mem_reg_194__3_ ( .D(n5547), .CK(clk), .QN(n2549) );
  DFF_X1 reg_mem_reg_194__2_ ( .D(n5546), .CK(clk), .QN(n2550) );
  DFF_X1 reg_mem_reg_194__1_ ( .D(n5545), .CK(clk), .QN(n2551) );
  DFF_X1 reg_mem_reg_194__0_ ( .D(n5544), .CK(clk), .QN(n2552) );
  DFF_X1 reg_mem_reg_195__7_ ( .D(n5543), .CK(clk), .QN(n2553) );
  DFF_X1 reg_mem_reg_195__6_ ( .D(n5542), .CK(clk), .QN(n2554) );
  DFF_X1 reg_mem_reg_195__5_ ( .D(n5541), .CK(clk), .QN(n2555) );
  DFF_X1 reg_mem_reg_195__4_ ( .D(n5540), .CK(clk), .QN(n2556) );
  DFF_X1 reg_mem_reg_195__3_ ( .D(n5539), .CK(clk), .QN(n2557) );
  DFF_X1 reg_mem_reg_195__2_ ( .D(n5538), .CK(clk), .QN(n2558) );
  DFF_X1 reg_mem_reg_195__1_ ( .D(n5537), .CK(clk), .QN(n2559) );
  DFF_X1 reg_mem_reg_195__0_ ( .D(n5536), .CK(clk), .QN(n2560) );
  DFF_X1 reg_mem_reg_196__7_ ( .D(n5535), .CK(clk), .Q(n[1040]), .QN(n2577) );
  DFF_X1 reg_mem_reg_196__6_ ( .D(n5534), .CK(clk), .Q(n[1039]), .QN(n2578) );
  DFF_X1 reg_mem_reg_196__5_ ( .D(n5533), .CK(clk), .Q(n[1038]), .QN(n2579) );
  DFF_X1 reg_mem_reg_196__4_ ( .D(n5532), .CK(clk), .Q(n[1037]), .QN(n2580) );
  DFF_X1 reg_mem_reg_196__3_ ( .D(n5531), .CK(clk), .Q(n[1036]), .QN(n2581) );
  DFF_X1 reg_mem_reg_196__2_ ( .D(n5530), .CK(clk), .Q(n[1035]), .QN(n2582) );
  DFF_X1 reg_mem_reg_196__1_ ( .D(n5529), .CK(clk), .Q(n[1034]), .QN(n2583) );
  DFF_X1 reg_mem_reg_196__0_ ( .D(n5528), .CK(clk), .Q(n[1033]), .QN(n2584) );
  DFF_X1 reg_mem_reg_197__7_ ( .D(n5527), .CK(clk), .Q(n[1032]), .QN(n2585) );
  DFF_X1 reg_mem_reg_197__6_ ( .D(n5526), .CK(clk), .Q(n[1031]), .QN(n2586) );
  DFF_X1 reg_mem_reg_197__5_ ( .D(n5525), .CK(clk), .Q(n[1030]), .QN(n2587) );
  DFF_X1 reg_mem_reg_197__4_ ( .D(n5524), .CK(clk), .Q(n[1029]), .QN(n2588) );
  DFF_X1 reg_mem_reg_197__3_ ( .D(n5523), .CK(clk), .Q(n[1028]), .QN(n2589) );
  DFF_X1 reg_mem_reg_197__2_ ( .D(n5522), .CK(clk), .Q(n[1027]), .QN(n2590) );
  DFF_X1 reg_mem_reg_197__1_ ( .D(n5521), .CK(clk), .Q(n[1026]), .QN(n2591) );
  DFF_X1 reg_mem_reg_197__0_ ( .D(n5520), .CK(clk), .Q(n[1025]), .QN(n2592) );
  DFF_X1 reg_mem_reg_198__7_ ( .D(n5519), .CK(clk), .QN(n2609) );
  DFF_X1 reg_mem_reg_198__6_ ( .D(n5518), .CK(clk), .QN(n2610) );
  DFF_X1 reg_mem_reg_198__5_ ( .D(n5517), .CK(clk), .QN(n2611) );
  DFF_X1 reg_mem_reg_198__4_ ( .D(n5516), .CK(clk), .QN(n2612) );
  DFF_X1 reg_mem_reg_198__3_ ( .D(n5515), .CK(clk), .QN(n2613) );
  DFF_X1 reg_mem_reg_198__2_ ( .D(n5514), .CK(clk), .QN(n2614) );
  DFF_X1 reg_mem_reg_198__1_ ( .D(n5513), .CK(clk), .QN(n2615) );
  DFF_X1 reg_mem_reg_198__0_ ( .D(n5512), .CK(clk), .QN(n2616) );
  DFF_X1 reg_mem_reg_199__7_ ( .D(n5511), .CK(clk), .QN(n2617) );
  DFF_X1 reg_mem_reg_199__6_ ( .D(n5510), .CK(clk), .QN(n2618) );
  DFF_X1 reg_mem_reg_199__5_ ( .D(n5509), .CK(clk), .QN(n2619) );
  DFF_X1 reg_mem_reg_199__4_ ( .D(n5508), .CK(clk), .QN(n2620) );
  DFF_X1 reg_mem_reg_199__3_ ( .D(n5507), .CK(clk), .QN(n2621) );
  DFF_X1 reg_mem_reg_199__2_ ( .D(n5506), .CK(clk), .QN(n2622) );
  DFF_X1 reg_mem_reg_199__1_ ( .D(n5505), .CK(clk), .QN(n2623) );
  DFF_X1 reg_mem_reg_199__0_ ( .D(n5504), .CK(clk), .QN(n2624) );
  DFF_X1 reg_mem_reg_200__7_ ( .D(n5503), .CK(clk), .Q(n[1008]), .QN(n2625) );
  DFF_X1 reg_mem_reg_200__6_ ( .D(n5502), .CK(clk), .Q(n[1007]), .QN(n2626) );
  DFF_X1 reg_mem_reg_200__5_ ( .D(n5501), .CK(clk), .Q(n[1006]), .QN(n2627) );
  DFF_X1 reg_mem_reg_200__4_ ( .D(n5500), .CK(clk), .Q(n[1005]), .QN(n2628) );
  DFF_X1 reg_mem_reg_200__3_ ( .D(n5499), .CK(clk), .Q(n[1004]), .QN(n2629) );
  DFF_X1 reg_mem_reg_200__2_ ( .D(n5498), .CK(clk), .Q(n[1003]), .QN(n2630) );
  DFF_X1 reg_mem_reg_200__1_ ( .D(n5497), .CK(clk), .Q(n[1002]), .QN(n2631) );
  DFF_X1 reg_mem_reg_200__0_ ( .D(n5496), .CK(clk), .Q(n[1001]), .QN(n2632) );
  DFF_X1 reg_mem_reg_201__7_ ( .D(n5495), .CK(clk), .Q(n[1000]), .QN(n2633) );
  DFF_X1 reg_mem_reg_201__6_ ( .D(n5494), .CK(clk), .Q(n[999]), .QN(n2634) );
  DFF_X1 reg_mem_reg_201__5_ ( .D(n5493), .CK(clk), .Q(n[998]), .QN(n2635) );
  DFF_X1 reg_mem_reg_201__4_ ( .D(n5492), .CK(clk), .Q(n[997]), .QN(n2636) );
  DFF_X1 reg_mem_reg_201__3_ ( .D(n5491), .CK(clk), .Q(n[996]), .QN(n2637) );
  DFF_X1 reg_mem_reg_201__2_ ( .D(n5490), .CK(clk), .Q(n[995]), .QN(n2638) );
  DFF_X1 reg_mem_reg_201__1_ ( .D(n5489), .CK(clk), .Q(n[994]), .QN(n2639) );
  DFF_X1 reg_mem_reg_201__0_ ( .D(n5488), .CK(clk), .Q(n[993]), .QN(n2640) );
  DFF_X1 reg_mem_reg_202__7_ ( .D(n5487), .CK(clk), .QN(n2641) );
  DFF_X1 reg_mem_reg_202__6_ ( .D(n5486), .CK(clk), .QN(n2642) );
  DFF_X1 reg_mem_reg_202__5_ ( .D(n5485), .CK(clk), .QN(n2643) );
  DFF_X1 reg_mem_reg_202__4_ ( .D(n5484), .CK(clk), .QN(n2644) );
  DFF_X1 reg_mem_reg_202__3_ ( .D(n5483), .CK(clk), .QN(n2645) );
  DFF_X1 reg_mem_reg_202__2_ ( .D(n5482), .CK(clk), .QN(n2646) );
  DFF_X1 reg_mem_reg_202__1_ ( .D(n5481), .CK(clk), .QN(n2647) );
  DFF_X1 reg_mem_reg_202__0_ ( .D(n5480), .CK(clk), .QN(n2648) );
  DFF_X1 reg_mem_reg_203__7_ ( .D(n5479), .CK(clk), .QN(n2649) );
  DFF_X1 reg_mem_reg_203__6_ ( .D(n5478), .CK(clk), .QN(n2650) );
  DFF_X1 reg_mem_reg_203__5_ ( .D(n5477), .CK(clk), .QN(n2651) );
  DFF_X1 reg_mem_reg_203__4_ ( .D(n5476), .CK(clk), .QN(n2652) );
  DFF_X1 reg_mem_reg_203__3_ ( .D(n5475), .CK(clk), .QN(n2653) );
  DFF_X1 reg_mem_reg_203__2_ ( .D(n5474), .CK(clk), .QN(n2654) );
  DFF_X1 reg_mem_reg_203__1_ ( .D(n5473), .CK(clk), .QN(n2655) );
  DFF_X1 reg_mem_reg_203__0_ ( .D(n5472), .CK(clk), .QN(n2656) );
  DFF_X1 reg_mem_reg_204__7_ ( .D(n5471), .CK(clk), .Q(n[976]), .QN(n2657) );
  DFF_X1 reg_mem_reg_204__6_ ( .D(n5470), .CK(clk), .Q(n[975]), .QN(n2658) );
  DFF_X1 reg_mem_reg_204__5_ ( .D(n5469), .CK(clk), .Q(n[974]), .QN(n2659) );
  DFF_X1 reg_mem_reg_204__4_ ( .D(n5468), .CK(clk), .Q(n[973]), .QN(n2660) );
  DFF_X1 reg_mem_reg_204__3_ ( .D(n5467), .CK(clk), .Q(n[972]), .QN(n2661) );
  DFF_X1 reg_mem_reg_204__2_ ( .D(n5466), .CK(clk), .Q(n[971]), .QN(n2662) );
  DFF_X1 reg_mem_reg_204__1_ ( .D(n5465), .CK(clk), .Q(n[970]), .QN(n2663) );
  DFF_X1 reg_mem_reg_204__0_ ( .D(n5464), .CK(clk), .Q(n[969]), .QN(n2664) );
  DFF_X1 reg_mem_reg_205__7_ ( .D(n5463), .CK(clk), .Q(n[968]), .QN(n2665) );
  DFF_X1 reg_mem_reg_205__6_ ( .D(n5462), .CK(clk), .Q(n[967]), .QN(n2666) );
  DFF_X1 reg_mem_reg_205__5_ ( .D(n5461), .CK(clk), .Q(n[966]), .QN(n2667) );
  DFF_X1 reg_mem_reg_205__4_ ( .D(n5460), .CK(clk), .Q(n[965]), .QN(n2668) );
  DFF_X1 reg_mem_reg_205__3_ ( .D(n5459), .CK(clk), .Q(n[964]), .QN(n2669) );
  DFF_X1 reg_mem_reg_205__2_ ( .D(n5458), .CK(clk), .Q(n[963]), .QN(n2670) );
  DFF_X1 reg_mem_reg_205__1_ ( .D(n5457), .CK(clk), .Q(n[962]), .QN(n2671) );
  DFF_X1 reg_mem_reg_205__0_ ( .D(n5456), .CK(clk), .Q(n[961]), .QN(n2672) );
  DFF_X1 reg_mem_reg_206__7_ ( .D(n5455), .CK(clk), .QN(n2673) );
  DFF_X1 reg_mem_reg_206__6_ ( .D(n5454), .CK(clk), .QN(n2674) );
  DFF_X1 reg_mem_reg_206__5_ ( .D(n5453), .CK(clk), .QN(n2675) );
  DFF_X1 reg_mem_reg_206__4_ ( .D(n5452), .CK(clk), .QN(n2676) );
  DFF_X1 reg_mem_reg_206__3_ ( .D(n5451), .CK(clk), .QN(n2677) );
  DFF_X1 reg_mem_reg_206__2_ ( .D(n5450), .CK(clk), .QN(n2678) );
  DFF_X1 reg_mem_reg_206__1_ ( .D(n5449), .CK(clk), .QN(n2679) );
  DFF_X1 reg_mem_reg_206__0_ ( .D(n5448), .CK(clk), .QN(n2680) );
  DFF_X1 reg_mem_reg_207__7_ ( .D(n5447), .CK(clk), .QN(n2681) );
  DFF_X1 reg_mem_reg_207__6_ ( .D(n5446), .CK(clk), .QN(n2682) );
  DFF_X1 reg_mem_reg_207__5_ ( .D(n5445), .CK(clk), .QN(n2683) );
  DFF_X1 reg_mem_reg_207__4_ ( .D(n5444), .CK(clk), .QN(n2684) );
  DFF_X1 reg_mem_reg_207__3_ ( .D(n5443), .CK(clk), .QN(n2685) );
  DFF_X1 reg_mem_reg_207__2_ ( .D(n5442), .CK(clk), .QN(n2686) );
  DFF_X1 reg_mem_reg_207__1_ ( .D(n5441), .CK(clk), .QN(n2687) );
  DFF_X1 reg_mem_reg_207__0_ ( .D(n5440), .CK(clk), .QN(n2688) );
  DFF_X1 reg_mem_reg_208__7_ ( .D(n5439), .CK(clk), .Q(n[944]), .QN(n2689) );
  DFF_X1 reg_mem_reg_208__6_ ( .D(n5438), .CK(clk), .Q(n[943]), .QN(n2690) );
  DFF_X1 reg_mem_reg_208__5_ ( .D(n5437), .CK(clk), .Q(n[942]), .QN(n2691) );
  DFF_X1 reg_mem_reg_208__4_ ( .D(n5436), .CK(clk), .Q(n[941]), .QN(n2692) );
  DFF_X1 reg_mem_reg_208__3_ ( .D(n5435), .CK(clk), .Q(n[940]), .QN(n2693) );
  DFF_X1 reg_mem_reg_208__2_ ( .D(n5434), .CK(clk), .Q(n[939]), .QN(n2694) );
  DFF_X1 reg_mem_reg_208__1_ ( .D(n5433), .CK(clk), .Q(n[938]), .QN(n2695) );
  DFF_X1 reg_mem_reg_208__0_ ( .D(n5432), .CK(clk), .Q(n[937]), .QN(n2696) );
  DFF_X1 reg_mem_reg_209__7_ ( .D(n5431), .CK(clk), .Q(n[936]), .QN(n2697) );
  DFF_X1 reg_mem_reg_209__6_ ( .D(n5430), .CK(clk), .Q(n[935]), .QN(n2698) );
  DFF_X1 reg_mem_reg_209__5_ ( .D(n5429), .CK(clk), .Q(n[934]), .QN(n2699) );
  DFF_X1 reg_mem_reg_209__4_ ( .D(n5428), .CK(clk), .Q(n[933]), .QN(n2700) );
  DFF_X1 reg_mem_reg_209__3_ ( .D(n5427), .CK(clk), .Q(n[932]), .QN(n2701) );
  DFF_X1 reg_mem_reg_209__2_ ( .D(n5426), .CK(clk), .Q(n[931]), .QN(n2702) );
  DFF_X1 reg_mem_reg_209__1_ ( .D(n5425), .CK(clk), .Q(n[930]), .QN(n2703) );
  DFF_X1 reg_mem_reg_209__0_ ( .D(n5424), .CK(clk), .Q(n[929]), .QN(n2704) );
  DFF_X1 reg_mem_reg_210__7_ ( .D(n5423), .CK(clk), .QN(n2705) );
  DFF_X1 reg_mem_reg_210__6_ ( .D(n5422), .CK(clk), .QN(n2706) );
  DFF_X1 reg_mem_reg_210__5_ ( .D(n5421), .CK(clk), .QN(n2707) );
  DFF_X1 reg_mem_reg_210__4_ ( .D(n5420), .CK(clk), .QN(n2708) );
  DFF_X1 reg_mem_reg_210__3_ ( .D(n5419), .CK(clk), .QN(n2709) );
  DFF_X1 reg_mem_reg_210__2_ ( .D(n5418), .CK(clk), .QN(n2710) );
  DFF_X1 reg_mem_reg_210__1_ ( .D(n5417), .CK(clk), .QN(n2711) );
  DFF_X1 reg_mem_reg_210__0_ ( .D(n5416), .CK(clk), .QN(n2712) );
  DFF_X1 reg_mem_reg_211__7_ ( .D(n5415), .CK(clk), .QN(n2713) );
  DFF_X1 reg_mem_reg_211__6_ ( .D(n5414), .CK(clk), .QN(n2714) );
  DFF_X1 reg_mem_reg_211__5_ ( .D(n5413), .CK(clk), .QN(n2715) );
  DFF_X1 reg_mem_reg_211__4_ ( .D(n5412), .CK(clk), .QN(n2716) );
  DFF_X1 reg_mem_reg_211__3_ ( .D(n5411), .CK(clk), .QN(n2717) );
  DFF_X1 reg_mem_reg_211__2_ ( .D(n5410), .CK(clk), .QN(n2718) );
  DFF_X1 reg_mem_reg_211__1_ ( .D(n5409), .CK(clk), .QN(n2719) );
  DFF_X1 reg_mem_reg_211__0_ ( .D(n5408), .CK(clk), .QN(n2720) );
  DFF_X1 reg_mem_reg_212__7_ ( .D(n5407), .CK(clk), .Q(n[912]), .QN(n2721) );
  DFF_X1 reg_mem_reg_212__6_ ( .D(n5406), .CK(clk), .Q(n[911]), .QN(n2722) );
  DFF_X1 reg_mem_reg_212__5_ ( .D(n5405), .CK(clk), .Q(n[910]), .QN(n2723) );
  DFF_X1 reg_mem_reg_212__4_ ( .D(n5404), .CK(clk), .Q(n[909]), .QN(n2724) );
  DFF_X1 reg_mem_reg_212__3_ ( .D(n5403), .CK(clk), .Q(n[908]), .QN(n2725) );
  DFF_X1 reg_mem_reg_212__2_ ( .D(n5402), .CK(clk), .Q(n[907]), .QN(n2726) );
  DFF_X1 reg_mem_reg_212__1_ ( .D(n5401), .CK(clk), .Q(n[906]), .QN(n2727) );
  DFF_X1 reg_mem_reg_212__0_ ( .D(n5400), .CK(clk), .Q(n[905]), .QN(n2728) );
  DFF_X1 reg_mem_reg_213__7_ ( .D(n5399), .CK(clk), .Q(n[904]), .QN(n2729) );
  DFF_X1 reg_mem_reg_213__6_ ( .D(n5398), .CK(clk), .Q(n[903]), .QN(n2730) );
  DFF_X1 reg_mem_reg_213__5_ ( .D(n5397), .CK(clk), .Q(n[902]), .QN(n2731) );
  DFF_X1 reg_mem_reg_213__4_ ( .D(n5396), .CK(clk), .Q(n[901]), .QN(n2732) );
  DFF_X1 reg_mem_reg_213__3_ ( .D(n5395), .CK(clk), .Q(n[900]), .QN(n2733) );
  DFF_X1 reg_mem_reg_213__2_ ( .D(n5394), .CK(clk), .Q(n[899]), .QN(n2734) );
  DFF_X1 reg_mem_reg_213__1_ ( .D(n5393), .CK(clk), .Q(n[898]), .QN(n2735) );
  DFF_X1 reg_mem_reg_213__0_ ( .D(n5392), .CK(clk), .Q(n[897]), .QN(n2736) );
  DFF_X1 reg_mem_reg_214__7_ ( .D(n5391), .CK(clk), .QN(n2737) );
  DFF_X1 reg_mem_reg_214__6_ ( .D(n5390), .CK(clk), .QN(n2738) );
  DFF_X1 reg_mem_reg_214__5_ ( .D(n5389), .CK(clk), .QN(n2739) );
  DFF_X1 reg_mem_reg_214__4_ ( .D(n5388), .CK(clk), .QN(n2740) );
  DFF_X1 reg_mem_reg_214__3_ ( .D(n5387), .CK(clk), .QN(n2741) );
  DFF_X1 reg_mem_reg_214__2_ ( .D(n5386), .CK(clk), .QN(n2742) );
  DFF_X1 reg_mem_reg_214__1_ ( .D(n5385), .CK(clk), .QN(n2743) );
  DFF_X1 reg_mem_reg_214__0_ ( .D(n5384), .CK(clk), .QN(n2744) );
  DFF_X1 reg_mem_reg_215__7_ ( .D(n5383), .CK(clk), .QN(n2745) );
  DFF_X1 reg_mem_reg_215__6_ ( .D(n5382), .CK(clk), .QN(n2746) );
  DFF_X1 reg_mem_reg_215__5_ ( .D(n5381), .CK(clk), .QN(n2747) );
  DFF_X1 reg_mem_reg_215__4_ ( .D(n5380), .CK(clk), .QN(n2748) );
  DFF_X1 reg_mem_reg_215__3_ ( .D(n5379), .CK(clk), .QN(n2749) );
  DFF_X1 reg_mem_reg_215__2_ ( .D(n5378), .CK(clk), .QN(n2750) );
  DFF_X1 reg_mem_reg_215__1_ ( .D(n5377), .CK(clk), .QN(n2751) );
  DFF_X1 reg_mem_reg_215__0_ ( .D(n5376), .CK(clk), .QN(n2752) );
  DFF_X1 reg_mem_reg_216__7_ ( .D(n5375), .CK(clk), .Q(n[880]), .QN(n2753) );
  DFF_X1 reg_mem_reg_216__6_ ( .D(n5374), .CK(clk), .Q(n[879]), .QN(n2754) );
  DFF_X1 reg_mem_reg_216__5_ ( .D(n5373), .CK(clk), .Q(n[878]), .QN(n2755) );
  DFF_X1 reg_mem_reg_216__4_ ( .D(n5372), .CK(clk), .Q(n[877]), .QN(n2756) );
  DFF_X1 reg_mem_reg_216__3_ ( .D(n5371), .CK(clk), .Q(n[876]), .QN(n2757) );
  DFF_X1 reg_mem_reg_216__2_ ( .D(n5370), .CK(clk), .Q(n[875]), .QN(n2758) );
  DFF_X1 reg_mem_reg_216__1_ ( .D(n5369), .CK(clk), .Q(n[874]), .QN(n2759) );
  DFF_X1 reg_mem_reg_216__0_ ( .D(n5368), .CK(clk), .Q(n[873]), .QN(n2760) );
  DFF_X1 reg_mem_reg_217__7_ ( .D(n5367), .CK(clk), .Q(n[872]), .QN(n2761) );
  DFF_X1 reg_mem_reg_217__6_ ( .D(n5366), .CK(clk), .Q(n[871]), .QN(n2762) );
  DFF_X1 reg_mem_reg_217__5_ ( .D(n5365), .CK(clk), .Q(n[870]), .QN(n2763) );
  DFF_X1 reg_mem_reg_217__4_ ( .D(n5364), .CK(clk), .Q(n[869]), .QN(n2764) );
  DFF_X1 reg_mem_reg_217__3_ ( .D(n5363), .CK(clk), .Q(n[868]), .QN(n2765) );
  DFF_X1 reg_mem_reg_217__2_ ( .D(n5362), .CK(clk), .Q(n[867]), .QN(n2766) );
  DFF_X1 reg_mem_reg_217__1_ ( .D(n5361), .CK(clk), .Q(n[866]), .QN(n2767) );
  DFF_X1 reg_mem_reg_217__0_ ( .D(n5360), .CK(clk), .Q(n[865]), .QN(n2768) );
  DFF_X1 reg_mem_reg_218__7_ ( .D(n5359), .CK(clk), .QN(n2769) );
  DFF_X1 reg_mem_reg_218__6_ ( .D(n5358), .CK(clk), .QN(n2770) );
  DFF_X1 reg_mem_reg_218__5_ ( .D(n5357), .CK(clk), .QN(n2771) );
  DFF_X1 reg_mem_reg_218__4_ ( .D(n5356), .CK(clk), .QN(n2772) );
  DFF_X1 reg_mem_reg_218__3_ ( .D(n5355), .CK(clk), .QN(n2773) );
  DFF_X1 reg_mem_reg_218__2_ ( .D(n5354), .CK(clk), .QN(n2774) );
  DFF_X1 reg_mem_reg_218__1_ ( .D(n5353), .CK(clk), .QN(n2775) );
  DFF_X1 reg_mem_reg_218__0_ ( .D(n5352), .CK(clk), .QN(n2776) );
  DFF_X1 reg_mem_reg_219__7_ ( .D(n5351), .CK(clk), .QN(n2777) );
  DFF_X1 reg_mem_reg_219__6_ ( .D(n5350), .CK(clk), .QN(n2778) );
  DFF_X1 reg_mem_reg_219__5_ ( .D(n5349), .CK(clk), .QN(n2779) );
  DFF_X1 reg_mem_reg_219__4_ ( .D(n5348), .CK(clk), .QN(n2780) );
  DFF_X1 reg_mem_reg_219__3_ ( .D(n5347), .CK(clk), .QN(n2781) );
  DFF_X1 reg_mem_reg_219__2_ ( .D(n5346), .CK(clk), .QN(n2782) );
  DFF_X1 reg_mem_reg_219__1_ ( .D(n5345), .CK(clk), .QN(n2783) );
  DFF_X1 reg_mem_reg_219__0_ ( .D(n5344), .CK(clk), .QN(n2784) );
  DFF_X1 reg_mem_reg_220__7_ ( .D(n5343), .CK(clk), .Q(n[848]), .QN(n2785) );
  DFF_X1 reg_mem_reg_220__6_ ( .D(n5342), .CK(clk), .Q(n[847]), .QN(n2786) );
  DFF_X1 reg_mem_reg_220__5_ ( .D(n5341), .CK(clk), .Q(n[846]), .QN(n2787) );
  DFF_X1 reg_mem_reg_220__4_ ( .D(n5340), .CK(clk), .Q(n[845]), .QN(n2788) );
  DFF_X1 reg_mem_reg_220__3_ ( .D(n5339), .CK(clk), .Q(n[844]), .QN(n2789) );
  DFF_X1 reg_mem_reg_220__2_ ( .D(n5338), .CK(clk), .Q(n[843]), .QN(n2790) );
  DFF_X1 reg_mem_reg_220__1_ ( .D(n5337), .CK(clk), .Q(n[842]), .QN(n2791) );
  DFF_X1 reg_mem_reg_220__0_ ( .D(n5336), .CK(clk), .Q(n[841]), .QN(n2792) );
  DFF_X1 reg_mem_reg_221__7_ ( .D(n5335), .CK(clk), .Q(n[840]), .QN(n2793) );
  DFF_X1 reg_mem_reg_221__6_ ( .D(n5334), .CK(clk), .Q(n[839]), .QN(n2794) );
  DFF_X1 reg_mem_reg_221__5_ ( .D(n5333), .CK(clk), .Q(n[838]), .QN(n2795) );
  DFF_X1 reg_mem_reg_221__4_ ( .D(n5332), .CK(clk), .Q(n[837]), .QN(n2796) );
  DFF_X1 reg_mem_reg_221__3_ ( .D(n5331), .CK(clk), .Q(n[836]), .QN(n2797) );
  DFF_X1 reg_mem_reg_221__2_ ( .D(n5330), .CK(clk), .Q(n[835]), .QN(n2798) );
  DFF_X1 reg_mem_reg_221__1_ ( .D(n5329), .CK(clk), .Q(n[834]), .QN(n2799) );
  DFF_X1 reg_mem_reg_221__0_ ( .D(n5328), .CK(clk), .Q(n[833]), .QN(n2800) );
  DFF_X1 reg_mem_reg_222__7_ ( .D(n5327), .CK(clk), .QN(n2801) );
  DFF_X1 reg_mem_reg_222__6_ ( .D(n5326), .CK(clk), .QN(n2802) );
  DFF_X1 reg_mem_reg_222__5_ ( .D(n5325), .CK(clk), .QN(n2803) );
  DFF_X1 reg_mem_reg_222__4_ ( .D(n5324), .CK(clk), .QN(n2804) );
  DFF_X1 reg_mem_reg_222__3_ ( .D(n5323), .CK(clk), .QN(n2805) );
  DFF_X1 reg_mem_reg_222__2_ ( .D(n5322), .CK(clk), .QN(n2806) );
  DFF_X1 reg_mem_reg_222__1_ ( .D(n5321), .CK(clk), .QN(n2807) );
  DFF_X1 reg_mem_reg_222__0_ ( .D(n5320), .CK(clk), .QN(n2808) );
  DFF_X1 reg_mem_reg_223__7_ ( .D(n5319), .CK(clk), .QN(n2809) );
  DFF_X1 reg_mem_reg_223__6_ ( .D(n5318), .CK(clk), .QN(n2810) );
  DFF_X1 reg_mem_reg_223__5_ ( .D(n5317), .CK(clk), .QN(n2811) );
  DFF_X1 reg_mem_reg_223__4_ ( .D(n5316), .CK(clk), .QN(n2812) );
  DFF_X1 reg_mem_reg_223__3_ ( .D(n5315), .CK(clk), .QN(n2813) );
  DFF_X1 reg_mem_reg_223__2_ ( .D(n5314), .CK(clk), .QN(n2814) );
  DFF_X1 reg_mem_reg_223__1_ ( .D(n5313), .CK(clk), .QN(n2815) );
  DFF_X1 reg_mem_reg_223__0_ ( .D(n5312), .CK(clk), .QN(n2816) );
  DFF_X1 reg_mem_reg_224__7_ ( .D(n5311), .CK(clk), .Q(n[816]), .QN(n2817) );
  DFF_X1 reg_mem_reg_224__6_ ( .D(n5310), .CK(clk), .Q(n[815]), .QN(n2818) );
  DFF_X1 reg_mem_reg_224__5_ ( .D(n5309), .CK(clk), .Q(n[814]), .QN(n2819) );
  DFF_X1 reg_mem_reg_224__4_ ( .D(n5308), .CK(clk), .Q(n[813]), .QN(n2820) );
  DFF_X1 reg_mem_reg_224__3_ ( .D(n5307), .CK(clk), .Q(n[812]), .QN(n2821) );
  DFF_X1 reg_mem_reg_224__2_ ( .D(n5306), .CK(clk), .Q(n[811]), .QN(n2822) );
  DFF_X1 reg_mem_reg_224__1_ ( .D(n5305), .CK(clk), .Q(n[810]), .QN(n2823) );
  DFF_X1 reg_mem_reg_224__0_ ( .D(n5304), .CK(clk), .Q(n[809]), .QN(n2824) );
  DFF_X1 reg_mem_reg_225__7_ ( .D(n5303), .CK(clk), .Q(n[808]), .QN(n2825) );
  DFF_X1 reg_mem_reg_225__6_ ( .D(n5302), .CK(clk), .Q(n[807]), .QN(n2826) );
  DFF_X1 reg_mem_reg_225__5_ ( .D(n5301), .CK(clk), .Q(n[806]), .QN(n2827) );
  DFF_X1 reg_mem_reg_225__4_ ( .D(n5300), .CK(clk), .Q(n[805]), .QN(n2828) );
  DFF_X1 reg_mem_reg_225__3_ ( .D(n5299), .CK(clk), .Q(n[804]), .QN(n2829) );
  DFF_X1 reg_mem_reg_225__2_ ( .D(n5298), .CK(clk), .Q(n[803]), .QN(n2830) );
  DFF_X1 reg_mem_reg_225__1_ ( .D(n5297), .CK(clk), .Q(n[802]), .QN(n2831) );
  DFF_X1 reg_mem_reg_225__0_ ( .D(n5296), .CK(clk), .Q(n[801]), .QN(n2832) );
  DFF_X1 reg_mem_reg_226__7_ ( .D(n5295), .CK(clk), .QN(n2833) );
  DFF_X1 reg_mem_reg_226__6_ ( .D(n5294), .CK(clk), .QN(n2834) );
  DFF_X1 reg_mem_reg_226__5_ ( .D(n5293), .CK(clk), .QN(n2835) );
  DFF_X1 reg_mem_reg_226__4_ ( .D(n5292), .CK(clk), .QN(n2836) );
  DFF_X1 reg_mem_reg_226__3_ ( .D(n5291), .CK(clk), .QN(n2837) );
  DFF_X1 reg_mem_reg_226__2_ ( .D(n5290), .CK(clk), .QN(n2838) );
  DFF_X1 reg_mem_reg_226__1_ ( .D(n5289), .CK(clk), .QN(n2839) );
  DFF_X1 reg_mem_reg_226__0_ ( .D(n5288), .CK(clk), .QN(n2840) );
  DFF_X1 reg_mem_reg_227__7_ ( .D(n5287), .CK(clk), .QN(n2841) );
  DFF_X1 reg_mem_reg_227__6_ ( .D(n5286), .CK(clk), .QN(n2842) );
  DFF_X1 reg_mem_reg_227__5_ ( .D(n5285), .CK(clk), .QN(n2843) );
  DFF_X1 reg_mem_reg_227__4_ ( .D(n5284), .CK(clk), .QN(n2844) );
  DFF_X1 reg_mem_reg_227__3_ ( .D(n5283), .CK(clk), .QN(n2845) );
  DFF_X1 reg_mem_reg_227__2_ ( .D(n5282), .CK(clk), .QN(n2846) );
  DFF_X1 reg_mem_reg_227__1_ ( .D(n5281), .CK(clk), .QN(n2847) );
  DFF_X1 reg_mem_reg_227__0_ ( .D(n5280), .CK(clk), .QN(n2848) );
  DFF_X1 reg_mem_reg_228__7_ ( .D(n5279), .CK(clk), .Q(n[784]), .QN(n2849) );
  DFF_X1 reg_mem_reg_228__6_ ( .D(n5278), .CK(clk), .Q(n[783]), .QN(n2850) );
  DFF_X1 reg_mem_reg_228__5_ ( .D(n5277), .CK(clk), .Q(n[782]), .QN(n2851) );
  DFF_X1 reg_mem_reg_228__4_ ( .D(n5276), .CK(clk), .Q(n[781]), .QN(n2852) );
  DFF_X1 reg_mem_reg_228__3_ ( .D(n5275), .CK(clk), .Q(n[780]), .QN(n2853) );
  DFF_X1 reg_mem_reg_228__2_ ( .D(n5274), .CK(clk), .Q(n[779]), .QN(n2854) );
  DFF_X1 reg_mem_reg_228__1_ ( .D(n5273), .CK(clk), .Q(n[778]), .QN(n2855) );
  DFF_X1 reg_mem_reg_228__0_ ( .D(n5272), .CK(clk), .Q(n[777]), .QN(n2856) );
  DFF_X1 reg_mem_reg_229__7_ ( .D(n5271), .CK(clk), .Q(n[776]), .QN(n2857) );
  DFF_X1 reg_mem_reg_229__6_ ( .D(n5270), .CK(clk), .Q(n[775]), .QN(n2858) );
  DFF_X1 reg_mem_reg_229__5_ ( .D(n5269), .CK(clk), .Q(n[774]), .QN(n2859) );
  DFF_X1 reg_mem_reg_229__4_ ( .D(n5268), .CK(clk), .Q(n[773]), .QN(n2860) );
  DFF_X1 reg_mem_reg_229__3_ ( .D(n5267), .CK(clk), .Q(n[772]), .QN(n2861) );
  DFF_X1 reg_mem_reg_229__2_ ( .D(n5266), .CK(clk), .Q(n[771]), .QN(n2862) );
  DFF_X1 reg_mem_reg_229__1_ ( .D(n5265), .CK(clk), .Q(n[770]), .QN(n2863) );
  DFF_X1 reg_mem_reg_229__0_ ( .D(n5264), .CK(clk), .Q(n[769]), .QN(n2864) );
  DFF_X1 reg_mem_reg_230__7_ ( .D(n5263), .CK(clk), .QN(n2865) );
  DFF_X1 reg_mem_reg_230__6_ ( .D(n5262), .CK(clk), .QN(n2866) );
  DFF_X1 reg_mem_reg_230__5_ ( .D(n5261), .CK(clk), .QN(n2867) );
  DFF_X1 reg_mem_reg_230__4_ ( .D(n5260), .CK(clk), .QN(n2868) );
  DFF_X1 reg_mem_reg_230__3_ ( .D(n5259), .CK(clk), .QN(n2869) );
  DFF_X1 reg_mem_reg_230__2_ ( .D(n5258), .CK(clk), .QN(n2870) );
  DFF_X1 reg_mem_reg_230__1_ ( .D(n5257), .CK(clk), .QN(n2871) );
  DFF_X1 reg_mem_reg_230__0_ ( .D(n5256), .CK(clk), .QN(n2872) );
  DFF_X1 reg_mem_reg_231__7_ ( .D(n5255), .CK(clk), .QN(n2873) );
  DFF_X1 reg_mem_reg_231__6_ ( .D(n5254), .CK(clk), .QN(n2874) );
  DFF_X1 reg_mem_reg_231__5_ ( .D(n5253), .CK(clk), .QN(n2875) );
  DFF_X1 reg_mem_reg_231__4_ ( .D(n5252), .CK(clk), .QN(n2876) );
  DFF_X1 reg_mem_reg_231__3_ ( .D(n5251), .CK(clk), .QN(n2877) );
  DFF_X1 reg_mem_reg_231__2_ ( .D(n5250), .CK(clk), .QN(n2878) );
  DFF_X1 reg_mem_reg_231__1_ ( .D(n5249), .CK(clk), .QN(n2879) );
  DFF_X1 reg_mem_reg_231__0_ ( .D(n5248), .CK(clk), .QN(n2880) );
  DFF_X1 reg_mem_reg_232__7_ ( .D(n5247), .CK(clk), .Q(n[752]), .QN(n2881) );
  DFF_X1 reg_mem_reg_232__6_ ( .D(n5246), .CK(clk), .Q(n[751]), .QN(n2882) );
  DFF_X1 reg_mem_reg_232__5_ ( .D(n5245), .CK(clk), .Q(n[750]), .QN(n2883) );
  DFF_X1 reg_mem_reg_232__4_ ( .D(n5244), .CK(clk), .Q(n[749]), .QN(n2884) );
  DFF_X1 reg_mem_reg_232__3_ ( .D(n5243), .CK(clk), .Q(n[748]), .QN(n2885) );
  DFF_X1 reg_mem_reg_232__2_ ( .D(n5242), .CK(clk), .Q(n[747]), .QN(n2886) );
  DFF_X1 reg_mem_reg_232__1_ ( .D(n5241), .CK(clk), .Q(n[746]), .QN(n2887) );
  DFF_X1 reg_mem_reg_232__0_ ( .D(n5240), .CK(clk), .Q(n[745]), .QN(n2888) );
  DFF_X1 reg_mem_reg_233__7_ ( .D(n5239), .CK(clk), .Q(n[744]), .QN(n2889) );
  DFF_X1 reg_mem_reg_233__6_ ( .D(n5238), .CK(clk), .Q(n[743]), .QN(n2890) );
  DFF_X1 reg_mem_reg_233__5_ ( .D(n5237), .CK(clk), .Q(n[742]), .QN(n2891) );
  DFF_X1 reg_mem_reg_233__4_ ( .D(n5236), .CK(clk), .Q(n[741]), .QN(n2892) );
  DFF_X1 reg_mem_reg_233__3_ ( .D(n5235), .CK(clk), .Q(n[740]), .QN(n2893) );
  DFF_X1 reg_mem_reg_233__2_ ( .D(n5234), .CK(clk), .Q(n[739]), .QN(n2894) );
  DFF_X1 reg_mem_reg_233__1_ ( .D(n5233), .CK(clk), .Q(n[738]), .QN(n2895) );
  DFF_X1 reg_mem_reg_233__0_ ( .D(n5232), .CK(clk), .Q(n[737]), .QN(n2896) );
  DFF_X1 reg_mem_reg_234__7_ ( .D(n5231), .CK(clk), .QN(n2897) );
  DFF_X1 reg_mem_reg_234__6_ ( .D(n5230), .CK(clk), .QN(n2898) );
  DFF_X1 reg_mem_reg_234__5_ ( .D(n5229), .CK(clk), .QN(n2899) );
  DFF_X1 reg_mem_reg_234__4_ ( .D(n5228), .CK(clk), .QN(n2900) );
  DFF_X1 reg_mem_reg_234__3_ ( .D(n5227), .CK(clk), .QN(n2901) );
  DFF_X1 reg_mem_reg_234__2_ ( .D(n5226), .CK(clk), .QN(n2902) );
  DFF_X1 reg_mem_reg_234__1_ ( .D(n5225), .CK(clk), .QN(n2903) );
  DFF_X1 reg_mem_reg_234__0_ ( .D(n5224), .CK(clk), .QN(n2904) );
  DFF_X1 reg_mem_reg_235__7_ ( .D(n5223), .CK(clk), .QN(n2905) );
  DFF_X1 reg_mem_reg_235__6_ ( .D(n5222), .CK(clk), .QN(n2906) );
  DFF_X1 reg_mem_reg_235__5_ ( .D(n5221), .CK(clk), .QN(n2907) );
  DFF_X1 reg_mem_reg_235__4_ ( .D(n5220), .CK(clk), .QN(n2908) );
  DFF_X1 reg_mem_reg_235__3_ ( .D(n5219), .CK(clk), .QN(n2909) );
  DFF_X1 reg_mem_reg_235__2_ ( .D(n5218), .CK(clk), .QN(n2910) );
  DFF_X1 reg_mem_reg_235__1_ ( .D(n5217), .CK(clk), .QN(n2911) );
  DFF_X1 reg_mem_reg_235__0_ ( .D(n5216), .CK(clk), .QN(n2912) );
  DFF_X1 reg_mem_reg_236__7_ ( .D(n5215), .CK(clk), .Q(n[720]), .QN(n2913) );
  DFF_X1 reg_mem_reg_236__6_ ( .D(n5214), .CK(clk), .Q(n[719]), .QN(n2914) );
  DFF_X1 reg_mem_reg_236__5_ ( .D(n5213), .CK(clk), .Q(n[718]), .QN(n2915) );
  DFF_X1 reg_mem_reg_236__4_ ( .D(n5212), .CK(clk), .Q(n[717]), .QN(n2916) );
  DFF_X1 reg_mem_reg_236__3_ ( .D(n5211), .CK(clk), .Q(n[716]), .QN(n2917) );
  DFF_X1 reg_mem_reg_236__2_ ( .D(n5210), .CK(clk), .Q(n[715]), .QN(n2918) );
  DFF_X1 reg_mem_reg_236__1_ ( .D(n5209), .CK(clk), .Q(n[714]), .QN(n2919) );
  DFF_X1 reg_mem_reg_236__0_ ( .D(n5208), .CK(clk), .Q(n[713]), .QN(n2920) );
  DFF_X1 reg_mem_reg_237__7_ ( .D(n5207), .CK(clk), .Q(n[712]), .QN(n2921) );
  DFF_X1 reg_mem_reg_237__6_ ( .D(n5206), .CK(clk), .Q(n[711]), .QN(n2922) );
  DFF_X1 reg_mem_reg_237__5_ ( .D(n5205), .CK(clk), .Q(n[710]), .QN(n2923) );
  DFF_X1 reg_mem_reg_237__4_ ( .D(n5204), .CK(clk), .Q(n[709]), .QN(n2924) );
  DFF_X1 reg_mem_reg_237__3_ ( .D(n5203), .CK(clk), .Q(n[708]), .QN(n2925) );
  DFF_X1 reg_mem_reg_237__2_ ( .D(n5202), .CK(clk), .Q(n[707]), .QN(n2926) );
  DFF_X1 reg_mem_reg_237__1_ ( .D(n5201), .CK(clk), .Q(n[706]), .QN(n2927) );
  DFF_X1 reg_mem_reg_237__0_ ( .D(n5200), .CK(clk), .Q(n[705]), .QN(n2928) );
  DFF_X1 reg_mem_reg_238__7_ ( .D(n5199), .CK(clk), .QN(n2929) );
  DFF_X1 reg_mem_reg_238__6_ ( .D(n5198), .CK(clk), .QN(n2930) );
  DFF_X1 reg_mem_reg_238__5_ ( .D(n5197), .CK(clk), .QN(n2931) );
  DFF_X1 reg_mem_reg_238__4_ ( .D(n5196), .CK(clk), .QN(n2932) );
  DFF_X1 reg_mem_reg_238__3_ ( .D(n5195), .CK(clk), .QN(n2933) );
  DFF_X1 reg_mem_reg_238__2_ ( .D(n5194), .CK(clk), .QN(n2934) );
  DFF_X1 reg_mem_reg_238__1_ ( .D(n5193), .CK(clk), .QN(n2935) );
  DFF_X1 reg_mem_reg_238__0_ ( .D(n5192), .CK(clk), .QN(n2936) );
  DFF_X1 reg_mem_reg_239__7_ ( .D(n5191), .CK(clk), .QN(n2937) );
  DFF_X1 reg_mem_reg_239__6_ ( .D(n5190), .CK(clk), .QN(n2938) );
  DFF_X1 reg_mem_reg_239__5_ ( .D(n5189), .CK(clk), .QN(n2939) );
  DFF_X1 reg_mem_reg_239__4_ ( .D(n5188), .CK(clk), .QN(n2940) );
  DFF_X1 reg_mem_reg_239__3_ ( .D(n5187), .CK(clk), .QN(n2941) );
  DFF_X1 reg_mem_reg_239__2_ ( .D(n5186), .CK(clk), .QN(n2942) );
  DFF_X1 reg_mem_reg_239__1_ ( .D(n5185), .CK(clk), .QN(n2943) );
  DFF_X1 reg_mem_reg_239__0_ ( .D(n5184), .CK(clk), .QN(n2944) );
  DFF_X1 reg_mem_reg_240__7_ ( .D(n5183), .CK(clk), .Q(n[688]), .QN(n2945) );
  DFF_X1 reg_mem_reg_240__6_ ( .D(n5182), .CK(clk), .Q(n[687]), .QN(n2946) );
  DFF_X1 reg_mem_reg_240__5_ ( .D(n5181), .CK(clk), .Q(n[686]), .QN(n2947) );
  DFF_X1 reg_mem_reg_240__4_ ( .D(n5180), .CK(clk), .Q(n[685]), .QN(n2948) );
  DFF_X1 reg_mem_reg_240__3_ ( .D(n5179), .CK(clk), .Q(n[684]), .QN(n2949) );
  DFF_X1 reg_mem_reg_240__2_ ( .D(n5178), .CK(clk), .Q(n[683]), .QN(n2950) );
  DFF_X1 reg_mem_reg_240__1_ ( .D(n5177), .CK(clk), .Q(n[682]), .QN(n2951) );
  DFF_X1 reg_mem_reg_240__0_ ( .D(n5176), .CK(clk), .Q(n[681]), .QN(n2952) );
  DFF_X1 reg_mem_reg_241__7_ ( .D(n5175), .CK(clk), .Q(n[680]), .QN(n2953) );
  DFF_X1 reg_mem_reg_241__6_ ( .D(n5174), .CK(clk), .Q(n[679]), .QN(n2954) );
  DFF_X1 reg_mem_reg_241__5_ ( .D(n5173), .CK(clk), .Q(n[678]), .QN(n2955) );
  DFF_X1 reg_mem_reg_241__4_ ( .D(n5172), .CK(clk), .Q(n[677]), .QN(n2956) );
  DFF_X1 reg_mem_reg_241__3_ ( .D(n5171), .CK(clk), .Q(n[676]), .QN(n2957) );
  DFF_X1 reg_mem_reg_241__2_ ( .D(n5170), .CK(clk), .Q(n[675]), .QN(n2958) );
  DFF_X1 reg_mem_reg_241__1_ ( .D(n5169), .CK(clk), .Q(n[674]), .QN(n2959) );
  DFF_X1 reg_mem_reg_241__0_ ( .D(n5168), .CK(clk), .Q(n[673]), .QN(n2960) );
  DFF_X1 reg_mem_reg_242__7_ ( .D(n5167), .CK(clk), .QN(n2961) );
  DFF_X1 reg_mem_reg_242__6_ ( .D(n5166), .CK(clk), .QN(n2962) );
  DFF_X1 reg_mem_reg_242__5_ ( .D(n5165), .CK(clk), .QN(n2963) );
  DFF_X1 reg_mem_reg_242__4_ ( .D(n5164), .CK(clk), .QN(n2964) );
  DFF_X1 reg_mem_reg_242__3_ ( .D(n5163), .CK(clk), .QN(n2965) );
  DFF_X1 reg_mem_reg_242__2_ ( .D(n5162), .CK(clk), .QN(n2966) );
  DFF_X1 reg_mem_reg_242__1_ ( .D(n5161), .CK(clk), .QN(n2967) );
  DFF_X1 reg_mem_reg_242__0_ ( .D(n5160), .CK(clk), .QN(n2968) );
  DFF_X1 reg_mem_reg_243__7_ ( .D(n5159), .CK(clk), .QN(n2969) );
  DFF_X1 reg_mem_reg_243__6_ ( .D(n5158), .CK(clk), .QN(n2970) );
  DFF_X1 reg_mem_reg_243__5_ ( .D(n5157), .CK(clk), .QN(n2971) );
  DFF_X1 reg_mem_reg_243__4_ ( .D(n5156), .CK(clk), .QN(n2972) );
  DFF_X1 reg_mem_reg_243__3_ ( .D(n5155), .CK(clk), .QN(n2973) );
  DFF_X1 reg_mem_reg_243__2_ ( .D(n5154), .CK(clk), .QN(n2974) );
  DFF_X1 reg_mem_reg_243__1_ ( .D(n5153), .CK(clk), .QN(n2975) );
  DFF_X1 reg_mem_reg_243__0_ ( .D(n5152), .CK(clk), .QN(n2976) );
  DFF_X1 reg_mem_reg_244__7_ ( .D(n5151), .CK(clk), .Q(n[656]), .QN(n2977) );
  DFF_X1 reg_mem_reg_244__6_ ( .D(n5150), .CK(clk), .Q(n[655]), .QN(n2978) );
  DFF_X1 reg_mem_reg_244__5_ ( .D(n5149), .CK(clk), .Q(n[654]), .QN(n2979) );
  DFF_X1 reg_mem_reg_244__4_ ( .D(n5148), .CK(clk), .Q(n[653]), .QN(n2980) );
  DFF_X1 reg_mem_reg_244__3_ ( .D(n5147), .CK(clk), .Q(n[652]), .QN(n2981) );
  DFF_X1 reg_mem_reg_244__2_ ( .D(n5146), .CK(clk), .Q(n[651]), .QN(n2982) );
  DFF_X1 reg_mem_reg_244__1_ ( .D(n5145), .CK(clk), .Q(n[650]), .QN(n2983) );
  DFF_X1 reg_mem_reg_244__0_ ( .D(n5144), .CK(clk), .Q(n[649]), .QN(n2984) );
  DFF_X1 reg_mem_reg_245__7_ ( .D(n5143), .CK(clk), .Q(n[648]), .QN(n2985) );
  DFF_X1 reg_mem_reg_245__6_ ( .D(n5142), .CK(clk), .Q(n[647]), .QN(n2986) );
  DFF_X1 reg_mem_reg_245__5_ ( .D(n5141), .CK(clk), .Q(n[646]), .QN(n2987) );
  DFF_X1 reg_mem_reg_245__4_ ( .D(n5140), .CK(clk), .Q(n[645]), .QN(n2988) );
  DFF_X1 reg_mem_reg_245__3_ ( .D(n5139), .CK(clk), .Q(n[644]), .QN(n2989) );
  DFF_X1 reg_mem_reg_245__2_ ( .D(n5138), .CK(clk), .Q(n[643]), .QN(n2990) );
  DFF_X1 reg_mem_reg_245__1_ ( .D(n5137), .CK(clk), .Q(n[642]), .QN(n2991) );
  DFF_X1 reg_mem_reg_245__0_ ( .D(n5136), .CK(clk), .Q(n[641]), .QN(n2992) );
  DFF_X1 reg_mem_reg_246__7_ ( .D(n5135), .CK(clk), .QN(n2993) );
  DFF_X1 reg_mem_reg_246__6_ ( .D(n5134), .CK(clk), .QN(n2994) );
  DFF_X1 reg_mem_reg_246__5_ ( .D(n5133), .CK(clk), .QN(n2995) );
  DFF_X1 reg_mem_reg_246__4_ ( .D(n5132), .CK(clk), .QN(n2996) );
  DFF_X1 reg_mem_reg_246__3_ ( .D(n5131), .CK(clk), .QN(n2997) );
  DFF_X1 reg_mem_reg_246__2_ ( .D(n5130), .CK(clk), .QN(n2998) );
  DFF_X1 reg_mem_reg_246__1_ ( .D(n5129), .CK(clk), .QN(n2999) );
  DFF_X1 reg_mem_reg_246__0_ ( .D(n5128), .CK(clk), .QN(n3000) );
  DFF_X1 reg_mem_reg_247__7_ ( .D(n5127), .CK(clk), .QN(n3001) );
  DFF_X1 reg_mem_reg_247__6_ ( .D(n5126), .CK(clk), .QN(n3002) );
  DFF_X1 reg_mem_reg_247__5_ ( .D(n5125), .CK(clk), .QN(n3003) );
  DFF_X1 reg_mem_reg_247__4_ ( .D(n5124), .CK(clk), .QN(n3004) );
  DFF_X1 reg_mem_reg_247__3_ ( .D(n5123), .CK(clk), .QN(n3005) );
  DFF_X1 reg_mem_reg_247__2_ ( .D(n5122), .CK(clk), .QN(n3006) );
  DFF_X1 reg_mem_reg_247__1_ ( .D(n5121), .CK(clk), .QN(n3007) );
  DFF_X1 reg_mem_reg_247__0_ ( .D(n5120), .CK(clk), .QN(n3008) );
  DFF_X1 reg_mem_reg_248__7_ ( .D(n5119), .CK(clk), .Q(n[624]), .QN(n3009) );
  DFF_X1 reg_mem_reg_248__6_ ( .D(n5118), .CK(clk), .Q(n[623]), .QN(n3010) );
  DFF_X1 reg_mem_reg_248__5_ ( .D(n5117), .CK(clk), .Q(n[622]), .QN(n3011) );
  DFF_X1 reg_mem_reg_248__4_ ( .D(n5116), .CK(clk), .Q(n[621]), .QN(n3012) );
  DFF_X1 reg_mem_reg_248__3_ ( .D(n5115), .CK(clk), .Q(n[620]), .QN(n3013) );
  DFF_X1 reg_mem_reg_248__2_ ( .D(n5114), .CK(clk), .Q(n[619]), .QN(n3014) );
  DFF_X1 reg_mem_reg_248__1_ ( .D(n5113), .CK(clk), .Q(n[618]), .QN(n3015) );
  DFF_X1 reg_mem_reg_248__0_ ( .D(n5112), .CK(clk), .Q(n[617]), .QN(n3016) );
  DFF_X1 reg_mem_reg_249__7_ ( .D(n5111), .CK(clk), .Q(n[616]), .QN(n3017) );
  DFF_X1 reg_mem_reg_249__6_ ( .D(n5110), .CK(clk), .Q(n[615]), .QN(n3018) );
  DFF_X1 reg_mem_reg_249__5_ ( .D(n5109), .CK(clk), .Q(n[614]), .QN(n3019) );
  DFF_X1 reg_mem_reg_249__4_ ( .D(n5108), .CK(clk), .Q(n[613]), .QN(n3020) );
  DFF_X1 reg_mem_reg_249__3_ ( .D(n5107), .CK(clk), .Q(n[612]), .QN(n3021) );
  DFF_X1 reg_mem_reg_249__2_ ( .D(n5106), .CK(clk), .Q(n[611]), .QN(n3022) );
  DFF_X1 reg_mem_reg_249__1_ ( .D(n5105), .CK(clk), .Q(n[610]), .QN(n3023) );
  DFF_X1 reg_mem_reg_249__0_ ( .D(n5104), .CK(clk), .Q(n[609]), .QN(n3024) );
  DFF_X1 reg_mem_reg_250__7_ ( .D(n5103), .CK(clk), .QN(n3025) );
  DFF_X1 reg_mem_reg_250__6_ ( .D(n5102), .CK(clk), .QN(n3026) );
  DFF_X1 reg_mem_reg_250__5_ ( .D(n5101), .CK(clk), .QN(n3027) );
  DFF_X1 reg_mem_reg_250__4_ ( .D(n5100), .CK(clk), .QN(n3028) );
  DFF_X1 reg_mem_reg_250__3_ ( .D(n5099), .CK(clk), .QN(n3029) );
  DFF_X1 reg_mem_reg_250__2_ ( .D(n5098), .CK(clk), .QN(n3030) );
  DFF_X1 reg_mem_reg_250__1_ ( .D(n5097), .CK(clk), .QN(n3031) );
  DFF_X1 reg_mem_reg_250__0_ ( .D(n5096), .CK(clk), .QN(n3032) );
  DFF_X1 reg_mem_reg_251__7_ ( .D(n5095), .CK(clk), .QN(n3033) );
  DFF_X1 reg_mem_reg_251__6_ ( .D(n5094), .CK(clk), .QN(n3034) );
  DFF_X1 reg_mem_reg_251__5_ ( .D(n5093), .CK(clk), .QN(n3035) );
  DFF_X1 reg_mem_reg_251__4_ ( .D(n5092), .CK(clk), .QN(n3036) );
  DFF_X1 reg_mem_reg_251__3_ ( .D(n5091), .CK(clk), .QN(n3037) );
  DFF_X1 reg_mem_reg_251__2_ ( .D(n5090), .CK(clk), .QN(n3038) );
  DFF_X1 reg_mem_reg_251__1_ ( .D(n5089), .CK(clk), .QN(n3039) );
  DFF_X1 reg_mem_reg_251__0_ ( .D(n5088), .CK(clk), .QN(n3040) );
  DFF_X1 reg_mem_reg_252__7_ ( .D(n5087), .CK(clk), .Q(n[592]), .QN(n3041) );
  DFF_X1 reg_mem_reg_252__6_ ( .D(n5086), .CK(clk), .Q(n[591]), .QN(n3042) );
  DFF_X1 reg_mem_reg_252__5_ ( .D(n5085), .CK(clk), .Q(n[590]), .QN(n3043) );
  DFF_X1 reg_mem_reg_252__4_ ( .D(n5084), .CK(clk), .Q(n[589]), .QN(n3044) );
  DFF_X1 reg_mem_reg_252__3_ ( .D(n5083), .CK(clk), .Q(n[588]), .QN(n3045) );
  DFF_X1 reg_mem_reg_252__2_ ( .D(n5082), .CK(clk), .Q(n[587]), .QN(n3046) );
  DFF_X1 reg_mem_reg_252__1_ ( .D(n5081), .CK(clk), .Q(n[586]), .QN(n3047) );
  DFF_X1 reg_mem_reg_252__0_ ( .D(n5080), .CK(clk), .Q(n[585]), .QN(n3048) );
  DFF_X1 reg_mem_reg_253__7_ ( .D(n5079), .CK(clk), .Q(n[584]), .QN(n3049) );
  DFF_X1 reg_mem_reg_253__6_ ( .D(n5078), .CK(clk), .Q(n[583]), .QN(n3050) );
  DFF_X1 reg_mem_reg_253__5_ ( .D(n5077), .CK(clk), .Q(n[582]), .QN(n3051) );
  DFF_X1 reg_mem_reg_253__4_ ( .D(n5076), .CK(clk), .Q(n[581]), .QN(n3052) );
  DFF_X1 reg_mem_reg_253__3_ ( .D(n5075), .CK(clk), .Q(n[580]), .QN(n3053) );
  DFF_X1 reg_mem_reg_253__2_ ( .D(n5074), .CK(clk), .Q(n[579]), .QN(n3054) );
  DFF_X1 reg_mem_reg_253__1_ ( .D(n5073), .CK(clk), .Q(n[578]), .QN(n3055) );
  DFF_X1 reg_mem_reg_253__0_ ( .D(n5072), .CK(clk), .Q(n[577]), .QN(n3056) );
  DFF_X1 reg_mem_reg_254__7_ ( .D(n5071), .CK(clk), .QN(n3057) );
  DFF_X1 reg_mem_reg_254__6_ ( .D(n5070), .CK(clk), .QN(n3058) );
  DFF_X1 reg_mem_reg_254__5_ ( .D(n5069), .CK(clk), .QN(n3059) );
  DFF_X1 reg_mem_reg_254__4_ ( .D(n5068), .CK(clk), .QN(n3060) );
  DFF_X1 reg_mem_reg_254__3_ ( .D(n5067), .CK(clk), .QN(n3061) );
  DFF_X1 reg_mem_reg_254__2_ ( .D(n5066), .CK(clk), .QN(n3062) );
  DFF_X1 reg_mem_reg_254__1_ ( .D(n5065), .CK(clk), .QN(n3063) );
  DFF_X1 reg_mem_reg_254__0_ ( .D(n5064), .CK(clk), .QN(n3064) );
  DFF_X1 reg_mem_reg_255__7_ ( .D(n5063), .CK(clk), .QN(n3065) );
  DFF_X1 reg_mem_reg_255__6_ ( .D(n5062), .CK(clk), .QN(n3066) );
  DFF_X1 reg_mem_reg_255__5_ ( .D(n5061), .CK(clk), .QN(n3067) );
  DFF_X1 reg_mem_reg_255__4_ ( .D(n5060), .CK(clk), .QN(n3068) );
  DFF_X1 reg_mem_reg_255__3_ ( .D(n5059), .CK(clk), .QN(n3069) );
  DFF_X1 reg_mem_reg_255__2_ ( .D(n5058), .CK(clk), .QN(n3070) );
  DFF_X1 reg_mem_reg_255__1_ ( .D(n5057), .CK(clk), .QN(n3071) );
  DFF_X1 reg_mem_reg_255__0_ ( .D(n5056), .CK(clk), .QN(n3072) );
  CLKBUF_X1 U2 ( .A(n3128), .Z(n3133) );
  CLKBUF_X1 U3 ( .A(n3128), .Z(n3132) );
  CLKBUF_X1 U4 ( .A(n3109), .Z(n3114) );
  CLKBUF_X1 U5 ( .A(n3109), .Z(n3115) );
  AND3_X1 U6 ( .A1(n3398), .A2(n3454), .A3(we_s), .ZN(n3352) );
  NOR2_X1 U7 ( .A1(n3232), .A2(addr_r[7]), .ZN(n3761) );
  NOR2_X1 U8 ( .A1(addr_r[6]), .A2(addr_r[7]), .ZN(n3804) );
  AND2_X1 U9 ( .A1(n3631), .A2(n3632), .ZN(n3351) );
  AND2_X1 U10 ( .A1(n3634), .A2(n3632), .ZN(n3354) );
  AND2_X1 U11 ( .A1(n3636), .A2(n3637), .ZN(n3356) );
  AND2_X1 U12 ( .A1(n3636), .A2(n3639), .ZN(n3358) );
  AND2_X1 U13 ( .A1(n3636), .A2(n3631), .ZN(n3360) );
  AND2_X1 U14 ( .A1(n3636), .A2(n3634), .ZN(n3362) );
  AND2_X1 U15 ( .A1(n3643), .A2(n3637), .ZN(n3364) );
  AND2_X1 U16 ( .A1(n3643), .A2(n3639), .ZN(n3366) );
  AND2_X1 U17 ( .A1(n3643), .A2(n3631), .ZN(n3368) );
  AND2_X1 U18 ( .A1(n3643), .A2(n3634), .ZN(n3370) );
  AND2_X1 U19 ( .A1(n3648), .A2(n3637), .ZN(n3372) );
  AND2_X1 U20 ( .A1(n3648), .A2(n3639), .ZN(n3374) );
  AND2_X1 U21 ( .A1(n3648), .A2(n3631), .ZN(n3376) );
  AND2_X1 U22 ( .A1(n3648), .A2(n3634), .ZN(n3378) );
  AND2_X1 U23 ( .A1(n3632), .A2(n3639), .ZN(n3383) );
  INV_X1 U24 ( .A(n3382), .ZN(n7132) );
  INV_X1 U25 ( .A(n3384), .ZN(n3295) );
  INV_X1 U26 ( .A(n3385), .ZN(n7243) );
  INV_X1 U27 ( .A(n3386), .ZN(n7114) );
  INV_X1 U28 ( .A(n3387), .ZN(n7179) );
  INV_X1 U29 ( .A(n3388), .ZN(n3279) );
  INV_X1 U30 ( .A(n3389), .ZN(n7227) );
  INV_X1 U31 ( .A(n3390), .ZN(n3343) );
  INV_X1 U32 ( .A(n3391), .ZN(n7163) );
  INV_X1 U33 ( .A(n3392), .ZN(n3263) );
  INV_X1 U34 ( .A(n3393), .ZN(n7211) );
  INV_X1 U35 ( .A(n3394), .ZN(n3327) );
  INV_X1 U36 ( .A(n3395), .ZN(n7147) );
  INV_X1 U37 ( .A(n3396), .ZN(n3247) );
  INV_X1 U38 ( .A(n3397), .ZN(n7195) );
  INV_X1 U39 ( .A(n3541), .ZN(n3303) );
  INV_X1 U40 ( .A(n3543), .ZN(n7123) );
  INV_X1 U41 ( .A(n3544), .ZN(n3286) );
  INV_X1 U42 ( .A(n3545), .ZN(n7234) );
  INV_X1 U43 ( .A(n3546), .ZN(n7105) );
  INV_X1 U44 ( .A(n3547), .ZN(n7170) );
  INV_X1 U45 ( .A(n3548), .ZN(n3270) );
  INV_X1 U46 ( .A(n3549), .ZN(n7218) );
  INV_X1 U47 ( .A(n3550), .ZN(n3334) );
  INV_X1 U48 ( .A(n3551), .ZN(n7154) );
  INV_X1 U49 ( .A(n3552), .ZN(n3254) );
  INV_X1 U50 ( .A(n3553), .ZN(n7202) );
  INV_X1 U51 ( .A(n3554), .ZN(n3318) );
  INV_X1 U52 ( .A(n3555), .ZN(n7138) );
  INV_X1 U53 ( .A(n3556), .ZN(n3238) );
  INV_X1 U54 ( .A(n3557), .ZN(n7186) );
  INV_X1 U55 ( .A(n3559), .ZN(n3302) );
  INV_X1 U56 ( .A(n3561), .ZN(n7122) );
  INV_X1 U57 ( .A(n3562), .ZN(n3285) );
  INV_X1 U58 ( .A(n3563), .ZN(n7233) );
  INV_X1 U59 ( .A(n3564), .ZN(n7104) );
  INV_X1 U60 ( .A(n3565), .ZN(n7169) );
  INV_X1 U61 ( .A(n3566), .ZN(n3269) );
  INV_X1 U62 ( .A(n3567), .ZN(n7217) );
  INV_X1 U63 ( .A(n3568), .ZN(n3333) );
  INV_X1 U64 ( .A(n3569), .ZN(n7153) );
  INV_X1 U65 ( .A(n3570), .ZN(n3253) );
  INV_X1 U66 ( .A(n3571), .ZN(n7201) );
  INV_X1 U67 ( .A(n3572), .ZN(n3317) );
  INV_X1 U68 ( .A(n3573), .ZN(n7137) );
  INV_X1 U69 ( .A(n3574), .ZN(n3237) );
  INV_X1 U70 ( .A(n3575), .ZN(n7185) );
  INV_X1 U71 ( .A(n3576), .ZN(n3301) );
  INV_X1 U72 ( .A(n3578), .ZN(n7121) );
  INV_X1 U73 ( .A(n3579), .ZN(n3284) );
  INV_X1 U74 ( .A(n3580), .ZN(n7232) );
  INV_X1 U75 ( .A(n3581), .ZN(n3348) );
  INV_X1 U76 ( .A(n3582), .ZN(n7168) );
  INV_X1 U77 ( .A(n3583), .ZN(n3268) );
  INV_X1 U78 ( .A(n3584), .ZN(n7216) );
  INV_X1 U79 ( .A(n3585), .ZN(n3332) );
  INV_X1 U80 ( .A(n3586), .ZN(n7152) );
  INV_X1 U81 ( .A(n3587), .ZN(n3252) );
  INV_X1 U82 ( .A(n3588), .ZN(n7200) );
  INV_X1 U83 ( .A(n3589), .ZN(n3316) );
  INV_X1 U84 ( .A(n3590), .ZN(n7136) );
  INV_X1 U85 ( .A(n3591), .ZN(n3236) );
  INV_X1 U86 ( .A(n3592), .ZN(n7184) );
  INV_X1 U87 ( .A(n3593), .ZN(n3300) );
  INV_X1 U88 ( .A(n3595), .ZN(n7120) );
  INV_X1 U89 ( .A(n3596), .ZN(n3283) );
  INV_X1 U90 ( .A(n3597), .ZN(n7231) );
  INV_X1 U91 ( .A(n3598), .ZN(n3347) );
  INV_X1 U92 ( .A(n3599), .ZN(n7167) );
  INV_X1 U93 ( .A(n3600), .ZN(n3267) );
  INV_X1 U94 ( .A(n3601), .ZN(n7215) );
  INV_X1 U95 ( .A(n3602), .ZN(n3331) );
  INV_X1 U96 ( .A(n3603), .ZN(n7151) );
  INV_X1 U97 ( .A(n3604), .ZN(n3251) );
  INV_X1 U98 ( .A(n3605), .ZN(n7199) );
  INV_X1 U99 ( .A(n3606), .ZN(n3315) );
  INV_X1 U100 ( .A(n3607), .ZN(n7135) );
  INV_X1 U101 ( .A(n3608), .ZN(n3235) );
  INV_X1 U102 ( .A(n3609), .ZN(n7183) );
  INV_X1 U103 ( .A(n3610), .ZN(n3299) );
  INV_X1 U104 ( .A(n3612), .ZN(n7119) );
  INV_X1 U105 ( .A(n3613), .ZN(n3282) );
  INV_X1 U106 ( .A(n3614), .ZN(n7230) );
  INV_X1 U107 ( .A(n3615), .ZN(n3346) );
  INV_X1 U108 ( .A(n3616), .ZN(n7166) );
  INV_X1 U109 ( .A(n3617), .ZN(n3266) );
  INV_X1 U110 ( .A(n3618), .ZN(n7214) );
  INV_X1 U111 ( .A(n3619), .ZN(n3330) );
  INV_X1 U112 ( .A(n3620), .ZN(n7150) );
  INV_X1 U113 ( .A(n3621), .ZN(n3250) );
  INV_X1 U114 ( .A(n3622), .ZN(n7198) );
  INV_X1 U115 ( .A(n3623), .ZN(n3314) );
  INV_X1 U116 ( .A(n3624), .ZN(n7134) );
  INV_X1 U117 ( .A(n3625), .ZN(n3234) );
  INV_X1 U118 ( .A(n3626), .ZN(n7182) );
  INV_X1 U119 ( .A(n3627), .ZN(n3298) );
  INV_X1 U120 ( .A(n3629), .ZN(n7118) );
  INV_X1 U121 ( .A(n3630), .ZN(n3281) );
  INV_X1 U122 ( .A(n3633), .ZN(n7229) );
  INV_X1 U123 ( .A(n3635), .ZN(n3345) );
  INV_X1 U124 ( .A(n3638), .ZN(n7165) );
  INV_X1 U125 ( .A(n3640), .ZN(n3265) );
  INV_X1 U126 ( .A(n3641), .ZN(n7213) );
  INV_X1 U127 ( .A(n3642), .ZN(n3329) );
  INV_X1 U128 ( .A(n3644), .ZN(n7149) );
  INV_X1 U129 ( .A(n3645), .ZN(n3249) );
  INV_X1 U130 ( .A(n3646), .ZN(n7197) );
  INV_X1 U131 ( .A(n3647), .ZN(n3313) );
  INV_X1 U132 ( .A(n3649), .ZN(n7133) );
  INV_X1 U133 ( .A(n3650), .ZN(n3233) );
  INV_X1 U134 ( .A(n3651), .ZN(n7181) );
  INV_X1 U135 ( .A(n3400), .ZN(n3311) );
  INV_X1 U136 ( .A(n3402), .ZN(n7131) );
  INV_X1 U137 ( .A(n3403), .ZN(n3294) );
  INV_X1 U138 ( .A(n3404), .ZN(n7242) );
  INV_X1 U139 ( .A(n3405), .ZN(n7113) );
  INV_X1 U140 ( .A(n3406), .ZN(n7178) );
  INV_X1 U141 ( .A(n3407), .ZN(n3278) );
  INV_X1 U142 ( .A(n3408), .ZN(n7226) );
  INV_X1 U143 ( .A(n3409), .ZN(n3342) );
  INV_X1 U144 ( .A(n3410), .ZN(n7162) );
  INV_X1 U145 ( .A(n3411), .ZN(n3262) );
  INV_X1 U146 ( .A(n3412), .ZN(n7210) );
  INV_X1 U147 ( .A(n3413), .ZN(n3326) );
  INV_X1 U148 ( .A(n3414), .ZN(n7146) );
  INV_X1 U149 ( .A(n3415), .ZN(n3246) );
  INV_X1 U150 ( .A(n3416), .ZN(n7194) );
  INV_X1 U151 ( .A(n3419), .ZN(n3310) );
  INV_X1 U152 ( .A(n3421), .ZN(n7130) );
  INV_X1 U153 ( .A(n3422), .ZN(n3293) );
  INV_X1 U154 ( .A(n3423), .ZN(n7241) );
  INV_X1 U155 ( .A(n3424), .ZN(n7112) );
  INV_X1 U156 ( .A(n3425), .ZN(n7177) );
  INV_X1 U157 ( .A(n3426), .ZN(n3277) );
  INV_X1 U158 ( .A(n3427), .ZN(n7225) );
  INV_X1 U159 ( .A(n3428), .ZN(n3341) );
  INV_X1 U160 ( .A(n3429), .ZN(n7161) );
  INV_X1 U161 ( .A(n3430), .ZN(n3261) );
  INV_X1 U162 ( .A(n3431), .ZN(n7209) );
  INV_X1 U163 ( .A(n3432), .ZN(n3325) );
  INV_X1 U164 ( .A(n3433), .ZN(n7145) );
  INV_X1 U165 ( .A(n3434), .ZN(n3245) );
  INV_X1 U166 ( .A(n3435), .ZN(n7193) );
  INV_X1 U167 ( .A(n3437), .ZN(n3309) );
  INV_X1 U168 ( .A(n3439), .ZN(n7129) );
  INV_X1 U169 ( .A(n3440), .ZN(n3292) );
  INV_X1 U170 ( .A(n3441), .ZN(n7240) );
  INV_X1 U171 ( .A(n3442), .ZN(n7111) );
  INV_X1 U172 ( .A(n3443), .ZN(n7176) );
  INV_X1 U173 ( .A(n3444), .ZN(n3276) );
  INV_X1 U174 ( .A(n3445), .ZN(n7224) );
  INV_X1 U175 ( .A(n3446), .ZN(n3340) );
  INV_X1 U176 ( .A(n3447), .ZN(n7160) );
  INV_X1 U177 ( .A(n3448), .ZN(n3260) );
  INV_X1 U178 ( .A(n3449), .ZN(n7208) );
  INV_X1 U179 ( .A(n3450), .ZN(n3324) );
  INV_X1 U180 ( .A(n3451), .ZN(n7144) );
  INV_X1 U181 ( .A(n3452), .ZN(n3244) );
  INV_X1 U182 ( .A(n3453), .ZN(n7192) );
  INV_X1 U183 ( .A(n3455), .ZN(n3308) );
  INV_X1 U184 ( .A(n3457), .ZN(n7128) );
  INV_X1 U185 ( .A(n3458), .ZN(n3291) );
  INV_X1 U186 ( .A(n3459), .ZN(n7239) );
  INV_X1 U187 ( .A(n3460), .ZN(n7110) );
  INV_X1 U188 ( .A(n3461), .ZN(n7175) );
  INV_X1 U189 ( .A(n3462), .ZN(n3275) );
  INV_X1 U190 ( .A(n3463), .ZN(n7223) );
  INV_X1 U191 ( .A(n3464), .ZN(n3339) );
  INV_X1 U192 ( .A(n3465), .ZN(n7159) );
  INV_X1 U193 ( .A(n3466), .ZN(n3259) );
  INV_X1 U194 ( .A(n3467), .ZN(n7207) );
  INV_X1 U195 ( .A(n3468), .ZN(n3323) );
  INV_X1 U196 ( .A(n3469), .ZN(n7143) );
  INV_X1 U197 ( .A(n3470), .ZN(n3243) );
  INV_X1 U198 ( .A(n3471), .ZN(n7191) );
  INV_X1 U199 ( .A(n3472), .ZN(n3307) );
  INV_X1 U200 ( .A(n3474), .ZN(n7127) );
  INV_X1 U201 ( .A(n3475), .ZN(n3290) );
  INV_X1 U202 ( .A(n3476), .ZN(n7238) );
  INV_X1 U203 ( .A(n3477), .ZN(n7109) );
  INV_X1 U204 ( .A(n3478), .ZN(n7174) );
  INV_X1 U205 ( .A(n3479), .ZN(n3274) );
  INV_X1 U206 ( .A(n3480), .ZN(n7222) );
  INV_X1 U207 ( .A(n3481), .ZN(n3338) );
  INV_X1 U208 ( .A(n3482), .ZN(n7158) );
  INV_X1 U209 ( .A(n3483), .ZN(n3258) );
  INV_X1 U210 ( .A(n3484), .ZN(n7206) );
  INV_X1 U211 ( .A(n3485), .ZN(n3322) );
  INV_X1 U212 ( .A(n3486), .ZN(n7142) );
  INV_X1 U213 ( .A(n3487), .ZN(n3242) );
  INV_X1 U214 ( .A(n3488), .ZN(n7190) );
  INV_X1 U215 ( .A(n3490), .ZN(n3306) );
  INV_X1 U216 ( .A(n3492), .ZN(n7126) );
  INV_X1 U217 ( .A(n3493), .ZN(n3289) );
  INV_X1 U218 ( .A(n3494), .ZN(n7237) );
  INV_X1 U219 ( .A(n3495), .ZN(n7108) );
  INV_X1 U220 ( .A(n3496), .ZN(n7173) );
  INV_X1 U221 ( .A(n3497), .ZN(n3273) );
  INV_X1 U222 ( .A(n3498), .ZN(n7221) );
  INV_X1 U223 ( .A(n3499), .ZN(n3337) );
  INV_X1 U224 ( .A(n3500), .ZN(n7157) );
  INV_X1 U225 ( .A(n3501), .ZN(n3257) );
  INV_X1 U226 ( .A(n3502), .ZN(n7205) );
  INV_X1 U227 ( .A(n3503), .ZN(n3321) );
  INV_X1 U228 ( .A(n3504), .ZN(n7141) );
  INV_X1 U229 ( .A(n3505), .ZN(n3241) );
  INV_X1 U230 ( .A(n3506), .ZN(n7189) );
  INV_X1 U231 ( .A(n3507), .ZN(n3305) );
  INV_X1 U232 ( .A(n3509), .ZN(n7125) );
  INV_X1 U233 ( .A(n3510), .ZN(n3288) );
  INV_X1 U234 ( .A(n3511), .ZN(n7236) );
  INV_X1 U235 ( .A(n3512), .ZN(n7107) );
  INV_X1 U236 ( .A(n3513), .ZN(n7172) );
  INV_X1 U237 ( .A(n3514), .ZN(n3272) );
  INV_X1 U238 ( .A(n3515), .ZN(n7220) );
  INV_X1 U239 ( .A(n3516), .ZN(n3336) );
  INV_X1 U240 ( .A(n3517), .ZN(n7156) );
  INV_X1 U241 ( .A(n3518), .ZN(n3256) );
  INV_X1 U242 ( .A(n3519), .ZN(n7204) );
  INV_X1 U243 ( .A(n3520), .ZN(n3320) );
  INV_X1 U244 ( .A(n3521), .ZN(n7140) );
  INV_X1 U245 ( .A(n3522), .ZN(n3240) );
  INV_X1 U246 ( .A(n3523), .ZN(n7188) );
  INV_X1 U247 ( .A(n3524), .ZN(n3304) );
  INV_X1 U248 ( .A(n3526), .ZN(n7124) );
  INV_X1 U249 ( .A(n3527), .ZN(n3287) );
  INV_X1 U250 ( .A(n3528), .ZN(n7235) );
  INV_X1 U251 ( .A(n3529), .ZN(n7106) );
  INV_X1 U252 ( .A(n3530), .ZN(n7171) );
  INV_X1 U253 ( .A(n3531), .ZN(n3271) );
  INV_X1 U254 ( .A(n3532), .ZN(n7219) );
  INV_X1 U255 ( .A(n3533), .ZN(n3335) );
  INV_X1 U256 ( .A(n3534), .ZN(n7155) );
  INV_X1 U257 ( .A(n3535), .ZN(n3255) );
  INV_X1 U258 ( .A(n3536), .ZN(n7203) );
  INV_X1 U259 ( .A(n3537), .ZN(n3319) );
  INV_X1 U260 ( .A(n3538), .ZN(n7139) );
  INV_X1 U261 ( .A(n3539), .ZN(n3239) );
  INV_X1 U262 ( .A(n3540), .ZN(n7187) );
  INV_X1 U263 ( .A(n3652), .ZN(n3297) );
  INV_X1 U264 ( .A(n3353), .ZN(n7244) );
  INV_X1 U265 ( .A(n3355), .ZN(n7115) );
  INV_X1 U266 ( .A(n3357), .ZN(n7180) );
  INV_X1 U267 ( .A(n3359), .ZN(n3280) );
  INV_X1 U268 ( .A(n3361), .ZN(n7228) );
  INV_X1 U269 ( .A(n3363), .ZN(n3344) );
  INV_X1 U270 ( .A(n3365), .ZN(n7164) );
  INV_X1 U271 ( .A(n3367), .ZN(n3264) );
  INV_X1 U272 ( .A(n3369), .ZN(n7212) );
  INV_X1 U273 ( .A(n3371), .ZN(n3328) );
  INV_X1 U274 ( .A(n3373), .ZN(n7148) );
  INV_X1 U275 ( .A(n3375), .ZN(n3248) );
  INV_X1 U276 ( .A(n3377), .ZN(n7196) );
  INV_X1 U277 ( .A(n3379), .ZN(n3312) );
  INV_X1 U278 ( .A(n3350), .ZN(n3296) );
  INV_X1 U279 ( .A(n3349), .ZN(n7117) );
  BUF_X1 U280 ( .A(n3172), .Z(n3176) );
  BUF_X1 U281 ( .A(n3172), .Z(n3179) );
  BUF_X1 U282 ( .A(n3172), .Z(n3178) );
  BUF_X1 U283 ( .A(n3172), .Z(n3177) );
  BUF_X1 U284 ( .A(n3153), .Z(n3160) );
  BUF_X1 U285 ( .A(n3153), .Z(n3159) );
  BUF_X1 U286 ( .A(n3153), .Z(n3158) );
  NAND2_X1 U287 ( .A1(n3381), .A2(n3383), .ZN(n3382) );
  NAND2_X1 U288 ( .A1(n3381), .A2(n3351), .ZN(n3384) );
  NAND2_X1 U289 ( .A1(n3381), .A2(n3354), .ZN(n3385) );
  NAND2_X1 U290 ( .A1(n3381), .A2(n3356), .ZN(n3386) );
  NAND2_X1 U291 ( .A1(n3381), .A2(n3358), .ZN(n3387) );
  NAND2_X1 U292 ( .A1(n3381), .A2(n3360), .ZN(n3388) );
  NAND2_X1 U293 ( .A1(n3381), .A2(n3362), .ZN(n3389) );
  NAND2_X1 U294 ( .A1(n3381), .A2(n3364), .ZN(n3390) );
  NAND2_X1 U295 ( .A1(n3381), .A2(n3366), .ZN(n3391) );
  NAND2_X1 U296 ( .A1(n3381), .A2(n3368), .ZN(n3392) );
  NAND2_X1 U297 ( .A1(n3381), .A2(n3370), .ZN(n3393) );
  NAND2_X1 U298 ( .A1(n3381), .A2(n3372), .ZN(n3394) );
  NAND2_X1 U299 ( .A1(n3381), .A2(n3374), .ZN(n3395) );
  NAND2_X1 U300 ( .A1(n3381), .A2(n3376), .ZN(n3396) );
  NAND2_X1 U301 ( .A1(n3381), .A2(n3378), .ZN(n3397) );
  NAND2_X1 U302 ( .A1(n3542), .A2(n3380), .ZN(n3541) );
  NAND2_X1 U303 ( .A1(n3542), .A2(n3383), .ZN(n3543) );
  NAND2_X1 U304 ( .A1(n3542), .A2(n3351), .ZN(n3544) );
  NAND2_X1 U305 ( .A1(n3542), .A2(n3354), .ZN(n3545) );
  NAND2_X1 U306 ( .A1(n3542), .A2(n3356), .ZN(n3546) );
  NAND2_X1 U307 ( .A1(n3542), .A2(n3358), .ZN(n3547) );
  NAND2_X1 U308 ( .A1(n3542), .A2(n3360), .ZN(n3548) );
  NAND2_X1 U309 ( .A1(n3542), .A2(n3362), .ZN(n3549) );
  NAND2_X1 U310 ( .A1(n3542), .A2(n3364), .ZN(n3550) );
  NAND2_X1 U311 ( .A1(n3542), .A2(n3366), .ZN(n3551) );
  NAND2_X1 U312 ( .A1(n3542), .A2(n3368), .ZN(n3552) );
  NAND2_X1 U313 ( .A1(n3542), .A2(n3370), .ZN(n3553) );
  NAND2_X1 U314 ( .A1(n3542), .A2(n3372), .ZN(n3554) );
  NAND2_X1 U315 ( .A1(n3542), .A2(n3374), .ZN(n3555) );
  NAND2_X1 U316 ( .A1(n3542), .A2(n3376), .ZN(n3556) );
  NAND2_X1 U317 ( .A1(n3542), .A2(n3378), .ZN(n3557) );
  NAND2_X1 U318 ( .A1(n3560), .A2(n3380), .ZN(n3559) );
  NAND2_X1 U319 ( .A1(n3560), .A2(n3383), .ZN(n3561) );
  NAND2_X1 U320 ( .A1(n3560), .A2(n3351), .ZN(n3562) );
  NAND2_X1 U321 ( .A1(n3560), .A2(n3354), .ZN(n3563) );
  NAND2_X1 U322 ( .A1(n3560), .A2(n3356), .ZN(n3564) );
  NAND2_X1 U323 ( .A1(n3560), .A2(n3358), .ZN(n3565) );
  NAND2_X1 U324 ( .A1(n3560), .A2(n3360), .ZN(n3566) );
  NAND2_X1 U325 ( .A1(n3560), .A2(n3362), .ZN(n3567) );
  NAND2_X1 U326 ( .A1(n3560), .A2(n3364), .ZN(n3568) );
  NAND2_X1 U327 ( .A1(n3560), .A2(n3366), .ZN(n3569) );
  NAND2_X1 U328 ( .A1(n3560), .A2(n3368), .ZN(n3570) );
  NAND2_X1 U329 ( .A1(n3560), .A2(n3370), .ZN(n3571) );
  NAND2_X1 U330 ( .A1(n3560), .A2(n3372), .ZN(n3572) );
  NAND2_X1 U331 ( .A1(n3560), .A2(n3374), .ZN(n3573) );
  NAND2_X1 U332 ( .A1(n3560), .A2(n3376), .ZN(n3574) );
  NAND2_X1 U333 ( .A1(n3560), .A2(n3378), .ZN(n3575) );
  NAND2_X1 U334 ( .A1(n3577), .A2(n3380), .ZN(n3576) );
  NAND2_X1 U335 ( .A1(n3577), .A2(n3383), .ZN(n3578) );
  NAND2_X1 U336 ( .A1(n3577), .A2(n3351), .ZN(n3579) );
  NAND2_X1 U337 ( .A1(n3577), .A2(n3354), .ZN(n3580) );
  NAND2_X1 U338 ( .A1(n3577), .A2(n3356), .ZN(n3581) );
  NAND2_X1 U339 ( .A1(n3577), .A2(n3358), .ZN(n3582) );
  NAND2_X1 U340 ( .A1(n3577), .A2(n3360), .ZN(n3583) );
  NAND2_X1 U341 ( .A1(n3577), .A2(n3362), .ZN(n3584) );
  NAND2_X1 U342 ( .A1(n3577), .A2(n3364), .ZN(n3585) );
  NAND2_X1 U343 ( .A1(n3577), .A2(n3366), .ZN(n3586) );
  NAND2_X1 U344 ( .A1(n3577), .A2(n3368), .ZN(n3587) );
  NAND2_X1 U345 ( .A1(n3577), .A2(n3370), .ZN(n3588) );
  NAND2_X1 U346 ( .A1(n3577), .A2(n3372), .ZN(n3589) );
  NAND2_X1 U347 ( .A1(n3577), .A2(n3374), .ZN(n3590) );
  NAND2_X1 U348 ( .A1(n3577), .A2(n3376), .ZN(n3591) );
  NAND2_X1 U349 ( .A1(n3577), .A2(n3378), .ZN(n3592) );
  NAND2_X1 U350 ( .A1(n3594), .A2(n3380), .ZN(n3593) );
  NAND2_X1 U351 ( .A1(n3594), .A2(n3383), .ZN(n3595) );
  NAND2_X1 U352 ( .A1(n3594), .A2(n3351), .ZN(n3596) );
  NAND2_X1 U353 ( .A1(n3594), .A2(n3354), .ZN(n3597) );
  NAND2_X1 U354 ( .A1(n3594), .A2(n3356), .ZN(n3598) );
  NAND2_X1 U355 ( .A1(n3594), .A2(n3358), .ZN(n3599) );
  NAND2_X1 U356 ( .A1(n3594), .A2(n3360), .ZN(n3600) );
  NAND2_X1 U357 ( .A1(n3594), .A2(n3362), .ZN(n3601) );
  NAND2_X1 U358 ( .A1(n3594), .A2(n3364), .ZN(n3602) );
  NAND2_X1 U359 ( .A1(n3594), .A2(n3366), .ZN(n3603) );
  NAND2_X1 U360 ( .A1(n3594), .A2(n3368), .ZN(n3604) );
  NAND2_X1 U361 ( .A1(n3594), .A2(n3370), .ZN(n3605) );
  NAND2_X1 U362 ( .A1(n3594), .A2(n3372), .ZN(n3606) );
  NAND2_X1 U363 ( .A1(n3594), .A2(n3374), .ZN(n3607) );
  NAND2_X1 U364 ( .A1(n3594), .A2(n3376), .ZN(n3608) );
  NAND2_X1 U365 ( .A1(n3594), .A2(n3378), .ZN(n3609) );
  NAND2_X1 U366 ( .A1(n3611), .A2(n3380), .ZN(n3610) );
  NAND2_X1 U367 ( .A1(n3611), .A2(n3383), .ZN(n3612) );
  NAND2_X1 U368 ( .A1(n3611), .A2(n3351), .ZN(n3613) );
  NAND2_X1 U369 ( .A1(n3611), .A2(n3354), .ZN(n3614) );
  NAND2_X1 U370 ( .A1(n3611), .A2(n3356), .ZN(n3615) );
  NAND2_X1 U371 ( .A1(n3611), .A2(n3358), .ZN(n3616) );
  NAND2_X1 U372 ( .A1(n3611), .A2(n3360), .ZN(n3617) );
  NAND2_X1 U373 ( .A1(n3611), .A2(n3362), .ZN(n3618) );
  NAND2_X1 U374 ( .A1(n3611), .A2(n3364), .ZN(n3619) );
  NAND2_X1 U375 ( .A1(n3611), .A2(n3366), .ZN(n3620) );
  NAND2_X1 U376 ( .A1(n3611), .A2(n3368), .ZN(n3621) );
  NAND2_X1 U377 ( .A1(n3611), .A2(n3370), .ZN(n3622) );
  NAND2_X1 U378 ( .A1(n3611), .A2(n3372), .ZN(n3623) );
  NAND2_X1 U379 ( .A1(n3611), .A2(n3374), .ZN(n3624) );
  NAND2_X1 U380 ( .A1(n3611), .A2(n3376), .ZN(n3625) );
  NAND2_X1 U381 ( .A1(n3611), .A2(n3378), .ZN(n3626) );
  NAND2_X1 U382 ( .A1(n3628), .A2(n3380), .ZN(n3627) );
  NAND2_X1 U383 ( .A1(n3628), .A2(n3383), .ZN(n3629) );
  NAND2_X1 U384 ( .A1(n3628), .A2(n3351), .ZN(n3630) );
  NAND2_X1 U385 ( .A1(n3628), .A2(n3354), .ZN(n3633) );
  NAND2_X1 U386 ( .A1(n3628), .A2(n3356), .ZN(n3635) );
  NAND2_X1 U387 ( .A1(n3628), .A2(n3358), .ZN(n3638) );
  NAND2_X1 U388 ( .A1(n3628), .A2(n3360), .ZN(n3640) );
  NAND2_X1 U389 ( .A1(n3628), .A2(n3362), .ZN(n3641) );
  NAND2_X1 U390 ( .A1(n3628), .A2(n3364), .ZN(n3642) );
  NAND2_X1 U391 ( .A1(n3628), .A2(n3366), .ZN(n3644) );
  NAND2_X1 U392 ( .A1(n3628), .A2(n3368), .ZN(n3645) );
  NAND2_X1 U393 ( .A1(n3628), .A2(n3370), .ZN(n3646) );
  NAND2_X1 U394 ( .A1(n3628), .A2(n3372), .ZN(n3647) );
  NAND2_X1 U395 ( .A1(n3628), .A2(n3374), .ZN(n3649) );
  NAND2_X1 U396 ( .A1(n3628), .A2(n3376), .ZN(n3650) );
  NAND2_X1 U397 ( .A1(n3628), .A2(n3378), .ZN(n3651) );
  NAND2_X1 U398 ( .A1(n3401), .A2(n3380), .ZN(n3400) );
  NAND2_X1 U399 ( .A1(n3401), .A2(n3383), .ZN(n3402) );
  NAND2_X1 U400 ( .A1(n3401), .A2(n3351), .ZN(n3403) );
  NAND2_X1 U401 ( .A1(n3401), .A2(n3354), .ZN(n3404) );
  NAND2_X1 U402 ( .A1(n3401), .A2(n3356), .ZN(n3405) );
  NAND2_X1 U403 ( .A1(n3401), .A2(n3358), .ZN(n3406) );
  NAND2_X1 U404 ( .A1(n3401), .A2(n3360), .ZN(n3407) );
  NAND2_X1 U405 ( .A1(n3401), .A2(n3362), .ZN(n3408) );
  NAND2_X1 U406 ( .A1(n3401), .A2(n3364), .ZN(n3409) );
  NAND2_X1 U407 ( .A1(n3401), .A2(n3366), .ZN(n3410) );
  NAND2_X1 U408 ( .A1(n3401), .A2(n3368), .ZN(n3411) );
  NAND2_X1 U409 ( .A1(n3401), .A2(n3370), .ZN(n3412) );
  NAND2_X1 U410 ( .A1(n3401), .A2(n3372), .ZN(n3413) );
  NAND2_X1 U411 ( .A1(n3401), .A2(n3374), .ZN(n3414) );
  NAND2_X1 U412 ( .A1(n3401), .A2(n3376), .ZN(n3415) );
  NAND2_X1 U413 ( .A1(n3401), .A2(n3378), .ZN(n3416) );
  NAND2_X1 U414 ( .A1(n3420), .A2(n3380), .ZN(n3419) );
  NAND2_X1 U415 ( .A1(n3420), .A2(n3383), .ZN(n3421) );
  NAND2_X1 U416 ( .A1(n3420), .A2(n3351), .ZN(n3422) );
  NAND2_X1 U417 ( .A1(n3420), .A2(n3354), .ZN(n3423) );
  NAND2_X1 U418 ( .A1(n3420), .A2(n3356), .ZN(n3424) );
  NAND2_X1 U419 ( .A1(n3420), .A2(n3358), .ZN(n3425) );
  NAND2_X1 U420 ( .A1(n3420), .A2(n3360), .ZN(n3426) );
  NAND2_X1 U421 ( .A1(n3420), .A2(n3362), .ZN(n3427) );
  NAND2_X1 U422 ( .A1(n3420), .A2(n3364), .ZN(n3428) );
  NAND2_X1 U423 ( .A1(n3420), .A2(n3366), .ZN(n3429) );
  NAND2_X1 U424 ( .A1(n3420), .A2(n3368), .ZN(n3430) );
  NAND2_X1 U425 ( .A1(n3420), .A2(n3370), .ZN(n3431) );
  NAND2_X1 U426 ( .A1(n3420), .A2(n3372), .ZN(n3432) );
  NAND2_X1 U427 ( .A1(n3420), .A2(n3374), .ZN(n3433) );
  NAND2_X1 U428 ( .A1(n3420), .A2(n3376), .ZN(n3434) );
  NAND2_X1 U429 ( .A1(n3420), .A2(n3378), .ZN(n3435) );
  NAND2_X1 U430 ( .A1(n3438), .A2(n3380), .ZN(n3437) );
  NAND2_X1 U431 ( .A1(n3438), .A2(n3383), .ZN(n3439) );
  NAND2_X1 U432 ( .A1(n3438), .A2(n3351), .ZN(n3440) );
  NAND2_X1 U433 ( .A1(n3438), .A2(n3354), .ZN(n3441) );
  NAND2_X1 U434 ( .A1(n3438), .A2(n3356), .ZN(n3442) );
  NAND2_X1 U435 ( .A1(n3438), .A2(n3358), .ZN(n3443) );
  NAND2_X1 U436 ( .A1(n3438), .A2(n3360), .ZN(n3444) );
  NAND2_X1 U437 ( .A1(n3438), .A2(n3362), .ZN(n3445) );
  NAND2_X1 U438 ( .A1(n3438), .A2(n3364), .ZN(n3446) );
  NAND2_X1 U439 ( .A1(n3438), .A2(n3366), .ZN(n3447) );
  NAND2_X1 U440 ( .A1(n3438), .A2(n3368), .ZN(n3448) );
  NAND2_X1 U441 ( .A1(n3438), .A2(n3370), .ZN(n3449) );
  NAND2_X1 U442 ( .A1(n3438), .A2(n3372), .ZN(n3450) );
  NAND2_X1 U443 ( .A1(n3438), .A2(n3374), .ZN(n3451) );
  NAND2_X1 U444 ( .A1(n3438), .A2(n3376), .ZN(n3452) );
  NAND2_X1 U445 ( .A1(n3438), .A2(n3378), .ZN(n3453) );
  NAND2_X1 U446 ( .A1(n3456), .A2(n3380), .ZN(n3455) );
  NAND2_X1 U447 ( .A1(n3456), .A2(n3383), .ZN(n3457) );
  NAND2_X1 U448 ( .A1(n3456), .A2(n3351), .ZN(n3458) );
  NAND2_X1 U449 ( .A1(n3456), .A2(n3354), .ZN(n3459) );
  NAND2_X1 U450 ( .A1(n3456), .A2(n3356), .ZN(n3460) );
  NAND2_X1 U451 ( .A1(n3456), .A2(n3358), .ZN(n3461) );
  NAND2_X1 U452 ( .A1(n3456), .A2(n3360), .ZN(n3462) );
  NAND2_X1 U453 ( .A1(n3456), .A2(n3362), .ZN(n3463) );
  NAND2_X1 U454 ( .A1(n3456), .A2(n3364), .ZN(n3464) );
  NAND2_X1 U455 ( .A1(n3456), .A2(n3366), .ZN(n3465) );
  NAND2_X1 U456 ( .A1(n3456), .A2(n3368), .ZN(n3466) );
  NAND2_X1 U457 ( .A1(n3456), .A2(n3370), .ZN(n3467) );
  NAND2_X1 U458 ( .A1(n3456), .A2(n3372), .ZN(n3468) );
  NAND2_X1 U459 ( .A1(n3456), .A2(n3374), .ZN(n3469) );
  NAND2_X1 U460 ( .A1(n3456), .A2(n3376), .ZN(n3470) );
  NAND2_X1 U461 ( .A1(n3456), .A2(n3378), .ZN(n3471) );
  NAND2_X1 U462 ( .A1(n3473), .A2(n3380), .ZN(n3472) );
  NAND2_X1 U463 ( .A1(n3473), .A2(n3383), .ZN(n3474) );
  NAND2_X1 U464 ( .A1(n3473), .A2(n3351), .ZN(n3475) );
  NAND2_X1 U465 ( .A1(n3473), .A2(n3354), .ZN(n3476) );
  NAND2_X1 U466 ( .A1(n3473), .A2(n3356), .ZN(n3477) );
  NAND2_X1 U467 ( .A1(n3473), .A2(n3358), .ZN(n3478) );
  NAND2_X1 U468 ( .A1(n3473), .A2(n3360), .ZN(n3479) );
  NAND2_X1 U469 ( .A1(n3473), .A2(n3362), .ZN(n3480) );
  NAND2_X1 U470 ( .A1(n3473), .A2(n3364), .ZN(n3481) );
  NAND2_X1 U471 ( .A1(n3473), .A2(n3366), .ZN(n3482) );
  NAND2_X1 U472 ( .A1(n3473), .A2(n3368), .ZN(n3483) );
  NAND2_X1 U473 ( .A1(n3473), .A2(n3370), .ZN(n3484) );
  NAND2_X1 U474 ( .A1(n3473), .A2(n3372), .ZN(n3485) );
  NAND2_X1 U475 ( .A1(n3473), .A2(n3374), .ZN(n3486) );
  NAND2_X1 U476 ( .A1(n3473), .A2(n3376), .ZN(n3487) );
  NAND2_X1 U477 ( .A1(n3473), .A2(n3378), .ZN(n3488) );
  NAND2_X1 U478 ( .A1(n3491), .A2(n3380), .ZN(n3490) );
  NAND2_X1 U479 ( .A1(n3491), .A2(n3383), .ZN(n3492) );
  NAND2_X1 U480 ( .A1(n3491), .A2(n3351), .ZN(n3493) );
  NAND2_X1 U481 ( .A1(n3491), .A2(n3354), .ZN(n3494) );
  NAND2_X1 U482 ( .A1(n3491), .A2(n3356), .ZN(n3495) );
  NAND2_X1 U483 ( .A1(n3491), .A2(n3358), .ZN(n3496) );
  NAND2_X1 U484 ( .A1(n3491), .A2(n3360), .ZN(n3497) );
  NAND2_X1 U485 ( .A1(n3491), .A2(n3362), .ZN(n3498) );
  NAND2_X1 U486 ( .A1(n3491), .A2(n3364), .ZN(n3499) );
  NAND2_X1 U487 ( .A1(n3491), .A2(n3366), .ZN(n3500) );
  NAND2_X1 U488 ( .A1(n3491), .A2(n3368), .ZN(n3501) );
  NAND2_X1 U489 ( .A1(n3491), .A2(n3370), .ZN(n3502) );
  NAND2_X1 U490 ( .A1(n3491), .A2(n3372), .ZN(n3503) );
  NAND2_X1 U491 ( .A1(n3491), .A2(n3374), .ZN(n3504) );
  NAND2_X1 U492 ( .A1(n3491), .A2(n3376), .ZN(n3505) );
  NAND2_X1 U493 ( .A1(n3491), .A2(n3378), .ZN(n3506) );
  NAND2_X1 U494 ( .A1(n3508), .A2(n3380), .ZN(n3507) );
  NAND2_X1 U495 ( .A1(n3508), .A2(n3383), .ZN(n3509) );
  NAND2_X1 U496 ( .A1(n3508), .A2(n3351), .ZN(n3510) );
  NAND2_X1 U497 ( .A1(n3508), .A2(n3354), .ZN(n3511) );
  NAND2_X1 U498 ( .A1(n3508), .A2(n3356), .ZN(n3512) );
  NAND2_X1 U499 ( .A1(n3508), .A2(n3358), .ZN(n3513) );
  NAND2_X1 U500 ( .A1(n3508), .A2(n3360), .ZN(n3514) );
  NAND2_X1 U501 ( .A1(n3508), .A2(n3362), .ZN(n3515) );
  NAND2_X1 U502 ( .A1(n3508), .A2(n3364), .ZN(n3516) );
  NAND2_X1 U503 ( .A1(n3508), .A2(n3366), .ZN(n3517) );
  NAND2_X1 U504 ( .A1(n3508), .A2(n3368), .ZN(n3518) );
  NAND2_X1 U505 ( .A1(n3508), .A2(n3370), .ZN(n3519) );
  NAND2_X1 U506 ( .A1(n3508), .A2(n3372), .ZN(n3520) );
  NAND2_X1 U507 ( .A1(n3508), .A2(n3374), .ZN(n3521) );
  NAND2_X1 U508 ( .A1(n3508), .A2(n3376), .ZN(n3522) );
  NAND2_X1 U509 ( .A1(n3508), .A2(n3378), .ZN(n3523) );
  NAND2_X1 U510 ( .A1(n3525), .A2(n3380), .ZN(n3524) );
  NAND2_X1 U511 ( .A1(n3525), .A2(n3383), .ZN(n3526) );
  NAND2_X1 U512 ( .A1(n3525), .A2(n3351), .ZN(n3527) );
  NAND2_X1 U513 ( .A1(n3525), .A2(n3354), .ZN(n3528) );
  NAND2_X1 U514 ( .A1(n3525), .A2(n3356), .ZN(n3529) );
  NAND2_X1 U515 ( .A1(n3525), .A2(n3358), .ZN(n3530) );
  NAND2_X1 U516 ( .A1(n3525), .A2(n3360), .ZN(n3531) );
  NAND2_X1 U517 ( .A1(n3525), .A2(n3362), .ZN(n3532) );
  NAND2_X1 U518 ( .A1(n3525), .A2(n3364), .ZN(n3533) );
  NAND2_X1 U519 ( .A1(n3525), .A2(n3366), .ZN(n3534) );
  NAND2_X1 U520 ( .A1(n3525), .A2(n3368), .ZN(n3535) );
  NAND2_X1 U521 ( .A1(n3525), .A2(n3370), .ZN(n3536) );
  NAND2_X1 U522 ( .A1(n3525), .A2(n3372), .ZN(n3537) );
  NAND2_X1 U523 ( .A1(n3525), .A2(n3374), .ZN(n3538) );
  NAND2_X1 U524 ( .A1(n3525), .A2(n3376), .ZN(n3539) );
  NAND2_X1 U525 ( .A1(n3525), .A2(n3378), .ZN(n3540) );
  NAND2_X1 U526 ( .A1(n3380), .A2(n3352), .ZN(n3652) );
  NAND2_X1 U527 ( .A1(n3354), .A2(n3352), .ZN(n3353) );
  NAND2_X1 U528 ( .A1(n3356), .A2(n3352), .ZN(n3355) );
  NAND2_X1 U529 ( .A1(n3358), .A2(n3352), .ZN(n3357) );
  NAND2_X1 U530 ( .A1(n3360), .A2(n3352), .ZN(n3359) );
  NAND2_X1 U531 ( .A1(n3362), .A2(n3352), .ZN(n3361) );
  NAND2_X1 U532 ( .A1(n3364), .A2(n3352), .ZN(n3363) );
  NAND2_X1 U533 ( .A1(n3366), .A2(n3352), .ZN(n3365) );
  NAND2_X1 U534 ( .A1(n3368), .A2(n3352), .ZN(n3367) );
  NAND2_X1 U535 ( .A1(n3370), .A2(n3352), .ZN(n3369) );
  NAND2_X1 U536 ( .A1(n3372), .A2(n3352), .ZN(n3371) );
  NAND2_X1 U537 ( .A1(n3374), .A2(n3352), .ZN(n3373) );
  NAND2_X1 U538 ( .A1(n3376), .A2(n3352), .ZN(n3375) );
  NAND2_X1 U539 ( .A1(n3378), .A2(n3352), .ZN(n3377) );
  NAND2_X1 U540 ( .A1(n3380), .A2(n3381), .ZN(n3379) );
  NAND2_X1 U541 ( .A1(n3351), .A2(n3352), .ZN(n3350) );
  NAND2_X1 U542 ( .A1(n3383), .A2(n3352), .ZN(n3349) );
  BUF_X1 U543 ( .A(n3666), .Z(n3227) );
  BUF_X1 U544 ( .A(n3679), .Z(n3152) );
  BUF_X1 U545 ( .A(n3684), .Z(n3151) );
  BUF_X1 U546 ( .A(n3209), .Z(n3213) );
  BUF_X1 U547 ( .A(n3209), .Z(n3216) );
  BUF_X1 U548 ( .A(n3209), .Z(n3215) );
  BUF_X1 U549 ( .A(n3209), .Z(n3214) );
  BUF_X1 U550 ( .A(n3670), .Z(n3207) );
  BUF_X1 U551 ( .A(n3675), .Z(n3170) );
  BUF_X1 U552 ( .A(n3670), .Z(n3206) );
  BUF_X1 U553 ( .A(n3675), .Z(n3169) );
  BUF_X1 U554 ( .A(n3670), .Z(n3205) );
  BUF_X1 U555 ( .A(n3675), .Z(n3168) );
  BUF_X1 U556 ( .A(n3667), .Z(n3225) );
  BUF_X1 U557 ( .A(n3689), .Z(n3150) );
  BUF_X1 U558 ( .A(n3673), .Z(n3172) );
  BUF_X1 U559 ( .A(n3671), .Z(n3190) );
  BUF_X1 U560 ( .A(n3676), .Z(n3153) );
  AND2_X1 U561 ( .A1(n3637), .A2(n3632), .ZN(n3380) );
  BUF_X1 U562 ( .A(n3137), .Z(n3142) );
  BUF_X1 U563 ( .A(n3121), .Z(n3124) );
  BUF_X1 U564 ( .A(n3100), .Z(n3103) );
  BUF_X1 U565 ( .A(n3082), .Z(n3088) );
  BUF_X1 U566 ( .A(n3073), .Z(n3079) );
  BUF_X1 U567 ( .A(n3137), .Z(n3141) );
  BUF_X1 U568 ( .A(n3119), .Z(n3123) );
  BUF_X1 U569 ( .A(n3100), .Z(n3104) );
  BUF_X1 U570 ( .A(n3093), .Z(n3097) );
  BUF_X1 U571 ( .A(n3082), .Z(n3089) );
  BUF_X1 U572 ( .A(n3073), .Z(n3080) );
  BUF_X1 U573 ( .A(n3106), .Z(n3105) );
  BUF_X1 U574 ( .A(n3091), .Z(n3098) );
  BUF_X1 U575 ( .A(n3128), .Z(n3134) );
  BUF_X1 U576 ( .A(n3118), .Z(n3122) );
  BUF_X1 U577 ( .A(n7254), .Z(n3106) );
  BUF_X1 U578 ( .A(n3091), .Z(n3099) );
  BUF_X1 U579 ( .A(n3104), .Z(n3107) );
  BUF_X1 U580 ( .A(n3111), .Z(n3116) );
  BUF_X1 U581 ( .A(n3101), .Z(n3108) );
  BUF_X1 U582 ( .A(n3128), .Z(n3131) );
  BUF_X1 U583 ( .A(n3139), .Z(n3140) );
  BUF_X1 U584 ( .A(n7255), .Z(n3110) );
  BUF_X1 U585 ( .A(n7255), .Z(n3111) );
  BUF_X1 U586 ( .A(n7252), .Z(n3084) );
  BUF_X1 U587 ( .A(n7251), .Z(n3075) );
  BUF_X1 U588 ( .A(n3119), .Z(n3120) );
  BUF_X1 U589 ( .A(n7258), .Z(n3139) );
  BUF_X1 U590 ( .A(n7256), .Z(n3121) );
  BUF_X1 U591 ( .A(n3092), .Z(n3093) );
  BUF_X1 U592 ( .A(n3109), .Z(n3112) );
  BUF_X1 U593 ( .A(n3100), .Z(n3101) );
  BUF_X1 U594 ( .A(n3092), .Z(n3094) );
  BUF_X1 U595 ( .A(n3082), .Z(n3085) );
  BUF_X1 U596 ( .A(n3073), .Z(n3076) );
  BUF_X1 U597 ( .A(n3137), .Z(n3144) );
  BUF_X1 U598 ( .A(n3118), .Z(n3126) );
  BUF_X1 U599 ( .A(n3109), .Z(n3113) );
  BUF_X1 U600 ( .A(n3094), .Z(n3095) );
  BUF_X1 U601 ( .A(n3082), .Z(n3086) );
  BUF_X1 U602 ( .A(n3073), .Z(n3077) );
  BUF_X1 U603 ( .A(n3137), .Z(n3143) );
  BUF_X1 U604 ( .A(n3129), .Z(n3135) );
  BUF_X1 U605 ( .A(n3118), .Z(n3125) );
  BUF_X1 U606 ( .A(n3100), .Z(n3102) );
  BUF_X1 U607 ( .A(n3094), .Z(n3096) );
  BUF_X1 U608 ( .A(n3082), .Z(n3087) );
  BUF_X1 U609 ( .A(n3073), .Z(n3078) );
  BUF_X1 U610 ( .A(n3110), .Z(n3117) );
  BUF_X1 U611 ( .A(n3084), .Z(n3090) );
  BUF_X1 U612 ( .A(n3075), .Z(n3081) );
  BUF_X1 U613 ( .A(n3137), .Z(n3145) );
  BUF_X1 U614 ( .A(n3129), .Z(n3136) );
  BUF_X1 U615 ( .A(n3118), .Z(n3127) );
  AND3_X1 U616 ( .A1(we_s), .A2(n3398), .A3(n3399), .ZN(n3381) );
  AND3_X1 U617 ( .A1(we_s), .A2(n3454), .A3(n3558), .ZN(n3577) );
  AND3_X1 U618 ( .A1(we_s), .A2(n3398), .A3(n3417), .ZN(n3611) );
  AND3_X1 U619 ( .A1(we_s), .A2(n3398), .A3(n3436), .ZN(n3628) );
  AND3_X1 U620 ( .A1(we_s), .A2(n3454), .A3(n3418), .ZN(n3438) );
  AND3_X1 U621 ( .A1(we_s), .A2(n3454), .A3(n3489), .ZN(n3508) );
  AND3_X1 U622 ( .A1(n3417), .A2(we_s), .A3(n3558), .ZN(n3542) );
  AND3_X1 U623 ( .A1(n3436), .A2(we_s), .A3(n3558), .ZN(n3560) );
  AND3_X1 U624 ( .A1(n3399), .A2(we_s), .A3(n3558), .ZN(n3594) );
  AND3_X1 U625 ( .A1(n3417), .A2(we_s), .A3(n3418), .ZN(n3401) );
  AND3_X1 U626 ( .A1(n3418), .A2(we_s), .A3(n3436), .ZN(n3420) );
  AND3_X1 U627 ( .A1(n3399), .A2(we_s), .A3(n3418), .ZN(n3456) );
  AND3_X1 U628 ( .A1(n3417), .A2(we_s), .A3(n3489), .ZN(n3473) );
  AND3_X1 U629 ( .A1(n3436), .A2(we_s), .A3(n3489), .ZN(n3491) );
  AND3_X1 U630 ( .A1(n3399), .A2(we_s), .A3(n3489), .ZN(n3525) );
  BUF_X1 U631 ( .A(n3698), .Z(n3149) );
  BUF_X1 U632 ( .A(n3708), .Z(n3147) );
  BUF_X1 U633 ( .A(n3713), .Z(n3146) );
  BUF_X1 U634 ( .A(n3703), .Z(n3148) );
  BUF_X1 U635 ( .A(n3668), .Z(n3209) );
  BUF_X1 U636 ( .A(n3672), .Z(n3181) );
  AND2_X1 U637 ( .A1(n5030), .A2(n3230), .ZN(n3689) );
  AND2_X1 U638 ( .A1(n5025), .A2(n3230), .ZN(n3684) );
  AND2_X1 U639 ( .A1(n5015), .A2(n3230), .ZN(n3666) );
  AND2_X1 U640 ( .A1(n5020), .A2(n3230), .ZN(n3679) );
  NAND2_X1 U641 ( .A1(n5055), .A2(n3228), .ZN(n3673) );
  NAND4_X1 U642 ( .A1(n4877), .A2(n4878), .A3(n4879), .A4(n4880), .ZN(
        data_r[0]) );
  OAI21_X1 U643 ( .B1(n5007), .B2(n5008), .A(n3804), .ZN(n4877) );
  OAI21_X1 U644 ( .B1(n4965), .B2(n4966), .A(n3761), .ZN(n4878) );
  OAI21_X1 U645 ( .B1(n4923), .B2(n4924), .A(n3718), .ZN(n4879) );
  NAND4_X1 U646 ( .A1(n4705), .A2(n4706), .A3(n4707), .A4(n4708), .ZN(
        data_r[1]) );
  OAI21_X1 U647 ( .B1(n4835), .B2(n4836), .A(n3804), .ZN(n4705) );
  OAI21_X1 U648 ( .B1(n4793), .B2(n4794), .A(n3761), .ZN(n4706) );
  OAI21_X1 U649 ( .B1(n4751), .B2(n4752), .A(n3718), .ZN(n4707) );
  NAND4_X1 U650 ( .A1(n4533), .A2(n4534), .A3(n4535), .A4(n4536), .ZN(
        data_r[2]) );
  OAI21_X1 U651 ( .B1(n4663), .B2(n4664), .A(n3804), .ZN(n4533) );
  OAI21_X1 U652 ( .B1(n4579), .B2(n4580), .A(n3718), .ZN(n4535) );
  OAI21_X1 U653 ( .B1(n4621), .B2(n4622), .A(n3761), .ZN(n4534) );
  NAND4_X1 U654 ( .A1(n4361), .A2(n4362), .A3(n4363), .A4(n4364), .ZN(
        data_r[3]) );
  OAI21_X1 U655 ( .B1(n4491), .B2(n4492), .A(n3804), .ZN(n4361) );
  OAI21_X1 U656 ( .B1(n4449), .B2(n4450), .A(n3761), .ZN(n4362) );
  OAI21_X1 U657 ( .B1(n4407), .B2(n4408), .A(n3718), .ZN(n4363) );
  NAND4_X1 U658 ( .A1(n4189), .A2(n4190), .A3(n4191), .A4(n4192), .ZN(
        data_r[4]) );
  OAI21_X1 U659 ( .B1(n4319), .B2(n4320), .A(n3804), .ZN(n4189) );
  OAI21_X1 U660 ( .B1(n4277), .B2(n4278), .A(n3761), .ZN(n4190) );
  OAI21_X1 U661 ( .B1(n4235), .B2(n4236), .A(n3718), .ZN(n4191) );
  NAND4_X1 U662 ( .A1(n4017), .A2(n4018), .A3(n4019), .A4(n4020), .ZN(
        data_r[5]) );
  OAI21_X1 U663 ( .B1(n4147), .B2(n4148), .A(n3804), .ZN(n4017) );
  OAI21_X1 U664 ( .B1(n4105), .B2(n4106), .A(n3761), .ZN(n4018) );
  OAI21_X1 U665 ( .B1(n4063), .B2(n4064), .A(n3718), .ZN(n4019) );
  NAND4_X1 U666 ( .A1(n3845), .A2(n3846), .A3(n3847), .A4(n3848), .ZN(
        data_r[6]) );
  OAI21_X1 U667 ( .B1(n3849), .B2(n3850), .A(n3659), .ZN(n3848) );
  OAI21_X1 U668 ( .B1(n3975), .B2(n3976), .A(n3804), .ZN(n3845) );
  OAI21_X1 U669 ( .B1(n3933), .B2(n3934), .A(n3761), .ZN(n3846) );
  NAND4_X1 U670 ( .A1(n3653), .A2(n3654), .A3(n3655), .A4(n3656), .ZN(
        data_r[7]) );
  OAI21_X1 U671 ( .B1(n3802), .B2(n3803), .A(n3804), .ZN(n3653) );
  OAI21_X1 U672 ( .B1(n3657), .B2(n3658), .A(n3659), .ZN(n3656) );
  OAI21_X1 U673 ( .B1(n3759), .B2(n3760), .A(n3761), .ZN(n3654) );
  AND2_X1 U674 ( .A1(n5052), .A2(n3228), .ZN(n3671) );
  AND2_X1 U675 ( .A1(n5054), .A2(n3228), .ZN(n3676) );
  NOR2_X1 U676 ( .A1(n7247), .A2(n7246), .ZN(n3632) );
  NOR2_X1 U677 ( .A1(n7116), .A2(n7245), .ZN(n3637) );
  NOR2_X1 U678 ( .A1(n7249), .A2(addr_w[7]), .ZN(n3418) );
  NOR2_X1 U679 ( .A1(n7249), .A2(n7250), .ZN(n3558) );
  INV_X1 U680 ( .A(addr_w[7]), .ZN(n7250) );
  BUF_X1 U681 ( .A(n3130), .Z(n3128) );
  BUF_X1 U682 ( .A(n3119), .Z(n3118) );
  BUF_X1 U683 ( .A(n3092), .Z(n3091) );
  BUF_X1 U684 ( .A(n3138), .Z(n3137) );
  BUF_X1 U685 ( .A(n3130), .Z(n3129) );
  BUF_X1 U686 ( .A(n7255), .Z(n3109) );
  BUF_X1 U687 ( .A(n7254), .Z(n3100) );
  BUF_X1 U688 ( .A(n3083), .Z(n3082) );
  BUF_X1 U689 ( .A(n3074), .Z(n3073) );
  NAND3_X1 U690 ( .A1(addr_r[0]), .A2(addr_r[2]), .A3(addr_r[1]), .ZN(n3667)
         );
  NAND3_X1 U691 ( .A1(addr_r[2]), .A2(n3228), .A3(addr_r[1]), .ZN(n3668) );
  INV_X1 U692 ( .A(addr_r[0]), .ZN(n3228) );
  INV_X1 U693 ( .A(addr_r[3]), .ZN(n3230) );
  NOR2_X1 U694 ( .A1(addr_r[1]), .A2(addr_r[2]), .ZN(n5052) );
  NAND2_X1 U695 ( .A1(n5055), .A2(addr_r[0]), .ZN(n3672) );
  NOR2_X1 U696 ( .A1(n3229), .A2(addr_r[1]), .ZN(n5054) );
  INV_X1 U697 ( .A(addr_r[2]), .ZN(n3229) );
  NAND4_X1 U698 ( .A1(n4925), .A2(n4926), .A3(n4927), .A4(n4928), .ZN(n4924)
         );
  OAI21_X1 U699 ( .B1(n4941), .B2(n4942), .A(n3689), .ZN(n4925) );
  OAI21_X1 U700 ( .B1(n4937), .B2(n4938), .A(n3151), .ZN(n4926) );
  OAI21_X1 U701 ( .B1(n4933), .B2(n4934), .A(n3152), .ZN(n4927) );
  NAND4_X1 U702 ( .A1(n4967), .A2(n4968), .A3(n4969), .A4(n4970), .ZN(n4966)
         );
  OAI21_X1 U703 ( .B1(n4983), .B2(n4984), .A(n3689), .ZN(n4967) );
  OAI21_X1 U704 ( .B1(n4979), .B2(n4980), .A(n3151), .ZN(n4968) );
  OAI21_X1 U705 ( .B1(n4975), .B2(n4976), .A(n3152), .ZN(n4969) );
  NAND4_X1 U706 ( .A1(n5009), .A2(n5010), .A3(n5011), .A4(n5012), .ZN(n5008)
         );
  OAI21_X1 U707 ( .B1(n5028), .B2(n5029), .A(n3689), .ZN(n5009) );
  OAI21_X1 U708 ( .B1(n5023), .B2(n5024), .A(n3151), .ZN(n5010) );
  OAI21_X1 U709 ( .B1(n5018), .B2(n5019), .A(n3152), .ZN(n5011) );
  NAND4_X1 U710 ( .A1(n4753), .A2(n4754), .A3(n4755), .A4(n4756), .ZN(n4752)
         );
  OAI21_X1 U711 ( .B1(n4769), .B2(n4770), .A(n3689), .ZN(n4753) );
  OAI21_X1 U712 ( .B1(n4765), .B2(n4766), .A(n3151), .ZN(n4754) );
  OAI21_X1 U713 ( .B1(n4761), .B2(n4762), .A(n3152), .ZN(n4755) );
  NAND4_X1 U714 ( .A1(n4795), .A2(n4796), .A3(n4797), .A4(n4798), .ZN(n4794)
         );
  OAI21_X1 U715 ( .B1(n4811), .B2(n4812), .A(n3689), .ZN(n4795) );
  OAI21_X1 U716 ( .B1(n4807), .B2(n4808), .A(n3151), .ZN(n4796) );
  OAI21_X1 U717 ( .B1(n4803), .B2(n4804), .A(n3152), .ZN(n4797) );
  NAND4_X1 U718 ( .A1(n4837), .A2(n4838), .A3(n4839), .A4(n4840), .ZN(n4836)
         );
  OAI21_X1 U719 ( .B1(n4853), .B2(n4854), .A(n3689), .ZN(n4837) );
  OAI21_X1 U720 ( .B1(n4849), .B2(n4850), .A(n3151), .ZN(n4838) );
  OAI21_X1 U721 ( .B1(n4845), .B2(n4846), .A(n3152), .ZN(n4839) );
  NAND4_X1 U722 ( .A1(n4623), .A2(n4624), .A3(n4625), .A4(n4626), .ZN(n4622)
         );
  OAI21_X1 U723 ( .B1(n4639), .B2(n4640), .A(n3689), .ZN(n4623) );
  OAI21_X1 U724 ( .B1(n4635), .B2(n4636), .A(n3684), .ZN(n4624) );
  OAI21_X1 U725 ( .B1(n4631), .B2(n4632), .A(n3679), .ZN(n4625) );
  NAND4_X1 U726 ( .A1(n4581), .A2(n4582), .A3(n4583), .A4(n4584), .ZN(n4580)
         );
  OAI21_X1 U727 ( .B1(n4597), .B2(n4598), .A(n3689), .ZN(n4581) );
  OAI21_X1 U728 ( .B1(n4593), .B2(n4594), .A(n3684), .ZN(n4582) );
  OAI21_X1 U729 ( .B1(n4589), .B2(n4590), .A(n3679), .ZN(n4583) );
  NAND4_X1 U730 ( .A1(n4665), .A2(n4666), .A3(n4667), .A4(n4668), .ZN(n4664)
         );
  OAI21_X1 U731 ( .B1(n4681), .B2(n4682), .A(n3689), .ZN(n4665) );
  OAI21_X1 U732 ( .B1(n4677), .B2(n4678), .A(n3684), .ZN(n4666) );
  OAI21_X1 U733 ( .B1(n4673), .B2(n4674), .A(n3679), .ZN(n4667) );
  NAND4_X1 U734 ( .A1(n4409), .A2(n4410), .A3(n4411), .A4(n4412), .ZN(n4408)
         );
  OAI21_X1 U735 ( .B1(n4425), .B2(n4426), .A(n3689), .ZN(n4409) );
  OAI21_X1 U736 ( .B1(n4421), .B2(n4422), .A(n3684), .ZN(n4410) );
  OAI21_X1 U737 ( .B1(n4417), .B2(n4418), .A(n3679), .ZN(n4411) );
  NAND4_X1 U738 ( .A1(n4451), .A2(n4452), .A3(n4453), .A4(n4454), .ZN(n4450)
         );
  OAI21_X1 U739 ( .B1(n4467), .B2(n4468), .A(n3689), .ZN(n4451) );
  OAI21_X1 U740 ( .B1(n4463), .B2(n4464), .A(n3684), .ZN(n4452) );
  OAI21_X1 U741 ( .B1(n4459), .B2(n4460), .A(n3679), .ZN(n4453) );
  NAND4_X1 U742 ( .A1(n4493), .A2(n4494), .A3(n4495), .A4(n4496), .ZN(n4492)
         );
  OAI21_X1 U743 ( .B1(n4509), .B2(n4510), .A(n3689), .ZN(n4493) );
  OAI21_X1 U744 ( .B1(n4505), .B2(n4506), .A(n3684), .ZN(n4494) );
  OAI21_X1 U745 ( .B1(n4501), .B2(n4502), .A(n3679), .ZN(n4495) );
  NAND4_X1 U746 ( .A1(n4237), .A2(n4238), .A3(n4239), .A4(n4240), .ZN(n4236)
         );
  OAI21_X1 U747 ( .B1(n4253), .B2(n4254), .A(n3689), .ZN(n4237) );
  OAI21_X1 U748 ( .B1(n4249), .B2(n4250), .A(n3684), .ZN(n4238) );
  OAI21_X1 U749 ( .B1(n4245), .B2(n4246), .A(n3679), .ZN(n4239) );
  NAND4_X1 U750 ( .A1(n4279), .A2(n4280), .A3(n4281), .A4(n4282), .ZN(n4278)
         );
  OAI21_X1 U751 ( .B1(n4295), .B2(n4296), .A(n3689), .ZN(n4279) );
  OAI21_X1 U752 ( .B1(n4291), .B2(n4292), .A(n3684), .ZN(n4280) );
  OAI21_X1 U753 ( .B1(n4287), .B2(n4288), .A(n3679), .ZN(n4281) );
  NAND4_X1 U754 ( .A1(n4321), .A2(n4322), .A3(n4323), .A4(n4324), .ZN(n4320)
         );
  OAI21_X1 U755 ( .B1(n4337), .B2(n4338), .A(n3689), .ZN(n4321) );
  OAI21_X1 U756 ( .B1(n4333), .B2(n4334), .A(n3684), .ZN(n4322) );
  OAI21_X1 U757 ( .B1(n4329), .B2(n4330), .A(n3679), .ZN(n4323) );
  NAND4_X1 U758 ( .A1(n4065), .A2(n4066), .A3(n4067), .A4(n4068), .ZN(n4064)
         );
  OAI21_X1 U759 ( .B1(n4081), .B2(n4082), .A(n3150), .ZN(n4065) );
  OAI21_X1 U760 ( .B1(n4077), .B2(n4078), .A(n3151), .ZN(n4066) );
  OAI21_X1 U761 ( .B1(n4073), .B2(n4074), .A(n3152), .ZN(n4067) );
  NAND4_X1 U762 ( .A1(n4107), .A2(n4108), .A3(n4109), .A4(n4110), .ZN(n4106)
         );
  OAI21_X1 U763 ( .B1(n4123), .B2(n4124), .A(n3150), .ZN(n4107) );
  OAI21_X1 U764 ( .B1(n4119), .B2(n4120), .A(n3684), .ZN(n4108) );
  OAI21_X1 U765 ( .B1(n4115), .B2(n4116), .A(n3679), .ZN(n4109) );
  NAND4_X1 U766 ( .A1(n4149), .A2(n4150), .A3(n4151), .A4(n4152), .ZN(n4148)
         );
  OAI21_X1 U767 ( .B1(n4165), .B2(n4166), .A(n3150), .ZN(n4149) );
  OAI21_X1 U768 ( .B1(n4161), .B2(n4162), .A(n3684), .ZN(n4150) );
  OAI21_X1 U769 ( .B1(n4157), .B2(n4158), .A(n3679), .ZN(n4151) );
  NAND4_X1 U770 ( .A1(n3935), .A2(n3936), .A3(n3937), .A4(n3938), .ZN(n3934)
         );
  OAI21_X1 U771 ( .B1(n3951), .B2(n3952), .A(n3150), .ZN(n3935) );
  OAI21_X1 U772 ( .B1(n3947), .B2(n3948), .A(n3684), .ZN(n3936) );
  OAI21_X1 U773 ( .B1(n3943), .B2(n3944), .A(n3679), .ZN(n3937) );
  NAND4_X1 U774 ( .A1(n3977), .A2(n3978), .A3(n3979), .A4(n3980), .ZN(n3976)
         );
  OAI21_X1 U775 ( .B1(n3993), .B2(n3994), .A(n3150), .ZN(n3977) );
  OAI21_X1 U776 ( .B1(n3989), .B2(n3990), .A(n3684), .ZN(n3978) );
  OAI21_X1 U777 ( .B1(n3985), .B2(n3986), .A(n3679), .ZN(n3979) );
  NAND4_X1 U778 ( .A1(n3851), .A2(n3852), .A3(n3853), .A4(n3854), .ZN(n3850)
         );
  OAI21_X1 U779 ( .B1(n3867), .B2(n3868), .A(n3150), .ZN(n3851) );
  OAI21_X1 U780 ( .B1(n3863), .B2(n3864), .A(n3151), .ZN(n3852) );
  OAI21_X1 U781 ( .B1(n3859), .B2(n3860), .A(n3152), .ZN(n3853) );
  NAND4_X1 U782 ( .A1(n3762), .A2(n3763), .A3(n3764), .A4(n3765), .ZN(n3760)
         );
  OAI21_X1 U783 ( .B1(n3778), .B2(n3779), .A(n3150), .ZN(n3762) );
  OAI21_X1 U784 ( .B1(n3774), .B2(n3775), .A(n3684), .ZN(n3763) );
  OAI21_X1 U785 ( .B1(n3770), .B2(n3771), .A(n3679), .ZN(n3764) );
  NAND4_X1 U786 ( .A1(n3660), .A2(n3661), .A3(n3662), .A4(n3663), .ZN(n3658)
         );
  OAI21_X1 U787 ( .B1(n3687), .B2(n3688), .A(n3150), .ZN(n3660) );
  OAI21_X1 U788 ( .B1(n3682), .B2(n3683), .A(n3151), .ZN(n3661) );
  OAI21_X1 U789 ( .B1(n3677), .B2(n3678), .A(n3152), .ZN(n3662) );
  NAND4_X1 U790 ( .A1(n3805), .A2(n3806), .A3(n3807), .A4(n3808), .ZN(n3803)
         );
  OAI21_X1 U791 ( .B1(n3821), .B2(n3822), .A(n3150), .ZN(n3805) );
  OAI21_X1 U792 ( .B1(n3817), .B2(n3818), .A(n3684), .ZN(n3806) );
  OAI21_X1 U793 ( .B1(n3813), .B2(n3814), .A(n3679), .ZN(n3807) );
  NOR2_X1 U794 ( .A1(addr_r[4]), .A2(addr_r[5]), .ZN(n5030) );
  NAND4_X1 U795 ( .A1(n4945), .A2(n4946), .A3(n4947), .A4(n4948), .ZN(n4923)
         );
  OAI21_X1 U796 ( .B1(n4961), .B2(n4962), .A(n3146), .ZN(n4945) );
  OAI21_X1 U797 ( .B1(n4957), .B2(n4958), .A(n3147), .ZN(n4946) );
  OAI21_X1 U798 ( .B1(n4953), .B2(n4954), .A(n3703), .ZN(n4947) );
  NAND4_X1 U799 ( .A1(n4987), .A2(n4988), .A3(n4989), .A4(n4990), .ZN(n4965)
         );
  OAI21_X1 U800 ( .B1(n5003), .B2(n5004), .A(n3146), .ZN(n4987) );
  OAI21_X1 U801 ( .B1(n4999), .B2(n5000), .A(n3147), .ZN(n4988) );
  OAI21_X1 U802 ( .B1(n4995), .B2(n4996), .A(n3703), .ZN(n4989) );
  NAND4_X1 U803 ( .A1(n5033), .A2(n5034), .A3(n5035), .A4(n5036), .ZN(n5007)
         );
  OAI21_X1 U804 ( .B1(n5049), .B2(n5050), .A(n3146), .ZN(n5033) );
  OAI21_X1 U805 ( .B1(n5045), .B2(n5046), .A(n3147), .ZN(n5034) );
  OAI21_X1 U806 ( .B1(n5041), .B2(n5042), .A(n3703), .ZN(n5035) );
  NAND4_X1 U807 ( .A1(n4773), .A2(n4774), .A3(n4775), .A4(n4776), .ZN(n4751)
         );
  OAI21_X1 U808 ( .B1(n4789), .B2(n4790), .A(n3146), .ZN(n4773) );
  OAI21_X1 U809 ( .B1(n4785), .B2(n4786), .A(n3147), .ZN(n4774) );
  OAI21_X1 U810 ( .B1(n4781), .B2(n4782), .A(n3703), .ZN(n4775) );
  NAND4_X1 U811 ( .A1(n4815), .A2(n4816), .A3(n4817), .A4(n4818), .ZN(n4793)
         );
  OAI21_X1 U812 ( .B1(n4831), .B2(n4832), .A(n3146), .ZN(n4815) );
  OAI21_X1 U813 ( .B1(n4827), .B2(n4828), .A(n3147), .ZN(n4816) );
  OAI21_X1 U814 ( .B1(n4823), .B2(n4824), .A(n3703), .ZN(n4817) );
  NAND4_X1 U815 ( .A1(n4857), .A2(n4858), .A3(n4859), .A4(n4860), .ZN(n4835)
         );
  OAI21_X1 U816 ( .B1(n4873), .B2(n4874), .A(n3146), .ZN(n4857) );
  OAI21_X1 U817 ( .B1(n4869), .B2(n4870), .A(n3147), .ZN(n4858) );
  OAI21_X1 U818 ( .B1(n4865), .B2(n4866), .A(n3703), .ZN(n4859) );
  NAND4_X1 U819 ( .A1(n4643), .A2(n4644), .A3(n4645), .A4(n4646), .ZN(n4621)
         );
  OAI21_X1 U820 ( .B1(n4659), .B2(n4660), .A(n3713), .ZN(n4643) );
  OAI21_X1 U821 ( .B1(n4655), .B2(n4656), .A(n3708), .ZN(n4644) );
  OAI21_X1 U822 ( .B1(n4651), .B2(n4652), .A(n3148), .ZN(n4645) );
  NAND4_X1 U823 ( .A1(n4601), .A2(n4602), .A3(n4603), .A4(n4604), .ZN(n4579)
         );
  OAI21_X1 U824 ( .B1(n4617), .B2(n4618), .A(n3713), .ZN(n4601) );
  OAI21_X1 U825 ( .B1(n4613), .B2(n4614), .A(n3708), .ZN(n4602) );
  OAI21_X1 U826 ( .B1(n4609), .B2(n4610), .A(n3148), .ZN(n4603) );
  NAND4_X1 U827 ( .A1(n4685), .A2(n4686), .A3(n4687), .A4(n4688), .ZN(n4663)
         );
  OAI21_X1 U828 ( .B1(n4701), .B2(n4702), .A(n3713), .ZN(n4685) );
  OAI21_X1 U829 ( .B1(n4697), .B2(n4698), .A(n3708), .ZN(n4686) );
  OAI21_X1 U830 ( .B1(n4693), .B2(n4694), .A(n3148), .ZN(n4687) );
  NAND4_X1 U831 ( .A1(n4257), .A2(n4258), .A3(n4259), .A4(n4260), .ZN(n4235)
         );
  OAI21_X1 U832 ( .B1(n4273), .B2(n4274), .A(n3713), .ZN(n4257) );
  OAI21_X1 U833 ( .B1(n4269), .B2(n4270), .A(n3708), .ZN(n4258) );
  OAI21_X1 U834 ( .B1(n4265), .B2(n4266), .A(n3148), .ZN(n4259) );
  NAND4_X1 U835 ( .A1(n4299), .A2(n4300), .A3(n4301), .A4(n4302), .ZN(n4277)
         );
  OAI21_X1 U836 ( .B1(n4315), .B2(n4316), .A(n3713), .ZN(n4299) );
  OAI21_X1 U837 ( .B1(n4311), .B2(n4312), .A(n3708), .ZN(n4300) );
  OAI21_X1 U838 ( .B1(n4307), .B2(n4308), .A(n3148), .ZN(n4301) );
  NAND4_X1 U839 ( .A1(n4085), .A2(n4086), .A3(n4087), .A4(n4088), .ZN(n4063)
         );
  OAI21_X1 U840 ( .B1(n4101), .B2(n4102), .A(n3146), .ZN(n4085) );
  OAI21_X1 U841 ( .B1(n4097), .B2(n4098), .A(n3147), .ZN(n4086) );
  OAI21_X1 U842 ( .B1(n4093), .B2(n4094), .A(n3703), .ZN(n4087) );
  NAND4_X1 U843 ( .A1(n4127), .A2(n4128), .A3(n4129), .A4(n4130), .ZN(n4105)
         );
  OAI21_X1 U844 ( .B1(n4143), .B2(n4144), .A(n3713), .ZN(n4127) );
  OAI21_X1 U845 ( .B1(n4139), .B2(n4140), .A(n3708), .ZN(n4128) );
  OAI21_X1 U846 ( .B1(n4135), .B2(n4136), .A(n3703), .ZN(n4129) );
  NAND4_X1 U847 ( .A1(n4169), .A2(n4170), .A3(n4171), .A4(n4172), .ZN(n4147)
         );
  OAI21_X1 U848 ( .B1(n4185), .B2(n4186), .A(n3713), .ZN(n4169) );
  OAI21_X1 U849 ( .B1(n4181), .B2(n4182), .A(n3708), .ZN(n4170) );
  OAI21_X1 U850 ( .B1(n4177), .B2(n4178), .A(n3703), .ZN(n4171) );
  NAND4_X1 U851 ( .A1(n3955), .A2(n3956), .A3(n3957), .A4(n3958), .ZN(n3933)
         );
  OAI21_X1 U852 ( .B1(n3971), .B2(n3972), .A(n3713), .ZN(n3955) );
  OAI21_X1 U853 ( .B1(n3967), .B2(n3968), .A(n3708), .ZN(n3956) );
  OAI21_X1 U854 ( .B1(n3963), .B2(n3964), .A(n3703), .ZN(n3957) );
  NAND4_X1 U855 ( .A1(n3997), .A2(n3998), .A3(n3999), .A4(n4000), .ZN(n3975)
         );
  OAI21_X1 U856 ( .B1(n4013), .B2(n4014), .A(n3713), .ZN(n3997) );
  OAI21_X1 U857 ( .B1(n4009), .B2(n4010), .A(n3708), .ZN(n3998) );
  OAI21_X1 U858 ( .B1(n4005), .B2(n4006), .A(n3703), .ZN(n3999) );
  NAND4_X1 U859 ( .A1(n4429), .A2(n4430), .A3(n4431), .A4(n4432), .ZN(n4407)
         );
  OAI21_X1 U860 ( .B1(n4445), .B2(n4446), .A(n3713), .ZN(n4429) );
  OAI21_X1 U861 ( .B1(n4441), .B2(n4442), .A(n3708), .ZN(n4430) );
  OAI21_X1 U862 ( .B1(n4437), .B2(n4438), .A(n3148), .ZN(n4431) );
  NAND4_X1 U863 ( .A1(n4471), .A2(n4472), .A3(n4473), .A4(n4474), .ZN(n4449)
         );
  OAI21_X1 U864 ( .B1(n4487), .B2(n4488), .A(n3713), .ZN(n4471) );
  OAI21_X1 U865 ( .B1(n4483), .B2(n4484), .A(n3708), .ZN(n4472) );
  OAI21_X1 U866 ( .B1(n4479), .B2(n4480), .A(n3148), .ZN(n4473) );
  NAND4_X1 U867 ( .A1(n4513), .A2(n4514), .A3(n4515), .A4(n4516), .ZN(n4491)
         );
  OAI21_X1 U868 ( .B1(n4529), .B2(n4530), .A(n3713), .ZN(n4513) );
  OAI21_X1 U869 ( .B1(n4525), .B2(n4526), .A(n3708), .ZN(n4514) );
  OAI21_X1 U870 ( .B1(n4521), .B2(n4522), .A(n3148), .ZN(n4515) );
  NAND4_X1 U871 ( .A1(n4341), .A2(n4342), .A3(n4343), .A4(n4344), .ZN(n4319)
         );
  OAI21_X1 U872 ( .B1(n4357), .B2(n4358), .A(n3713), .ZN(n4341) );
  OAI21_X1 U873 ( .B1(n4353), .B2(n4354), .A(n3708), .ZN(n4342) );
  OAI21_X1 U874 ( .B1(n4349), .B2(n4350), .A(n3148), .ZN(n4343) );
  NAND4_X1 U875 ( .A1(n3871), .A2(n3872), .A3(n3873), .A4(n3874), .ZN(n3849)
         );
  OAI21_X1 U876 ( .B1(n3887), .B2(n3888), .A(n3146), .ZN(n3871) );
  OAI21_X1 U877 ( .B1(n3883), .B2(n3884), .A(n3147), .ZN(n3872) );
  OAI21_X1 U878 ( .B1(n3879), .B2(n3880), .A(n3703), .ZN(n3873) );
  NAND4_X1 U879 ( .A1(n3782), .A2(n3783), .A3(n3784), .A4(n3785), .ZN(n3759)
         );
  OAI21_X1 U880 ( .B1(n3798), .B2(n3799), .A(n3713), .ZN(n3782) );
  OAI21_X1 U881 ( .B1(n3794), .B2(n3795), .A(n3708), .ZN(n3783) );
  OAI21_X1 U882 ( .B1(n3790), .B2(n3791), .A(n3703), .ZN(n3784) );
  NAND4_X1 U883 ( .A1(n3692), .A2(n3693), .A3(n3694), .A4(n3695), .ZN(n3657)
         );
  OAI21_X1 U884 ( .B1(n3711), .B2(n3712), .A(n3146), .ZN(n3692) );
  OAI21_X1 U885 ( .B1(n3706), .B2(n3707), .A(n3147), .ZN(n3693) );
  OAI21_X1 U886 ( .B1(n3701), .B2(n3702), .A(n3703), .ZN(n3694) );
  NAND4_X1 U887 ( .A1(n3825), .A2(n3826), .A3(n3827), .A4(n3828), .ZN(n3802)
         );
  OAI21_X1 U888 ( .B1(n3841), .B2(n3842), .A(n3713), .ZN(n3825) );
  OAI21_X1 U889 ( .B1(n3837), .B2(n3838), .A(n3708), .ZN(n3826) );
  OAI21_X1 U890 ( .B1(n3833), .B2(n3834), .A(n3703), .ZN(n3827) );
  INV_X1 U891 ( .A(addr_r[4]), .ZN(n3231) );
  OAI21_X1 U892 ( .B1(n4881), .B2(n4882), .A(n3659), .ZN(n4880) );
  NAND4_X1 U893 ( .A1(n4903), .A2(n4904), .A3(n4905), .A4(n4906), .ZN(n4881)
         );
  NAND4_X1 U894 ( .A1(n4883), .A2(n4884), .A3(n4885), .A4(n4886), .ZN(n4882)
         );
  OAI21_X1 U895 ( .B1(n4919), .B2(n4920), .A(n3146), .ZN(n4903) );
  OAI21_X1 U896 ( .B1(n4709), .B2(n4710), .A(n3659), .ZN(n4708) );
  NAND4_X1 U897 ( .A1(n4731), .A2(n4732), .A3(n4733), .A4(n4734), .ZN(n4709)
         );
  NAND4_X1 U898 ( .A1(n4711), .A2(n4712), .A3(n4713), .A4(n4714), .ZN(n4710)
         );
  OAI21_X1 U899 ( .B1(n4747), .B2(n4748), .A(n3146), .ZN(n4731) );
  OAI21_X1 U900 ( .B1(n4537), .B2(n4538), .A(n3659), .ZN(n4536) );
  NAND4_X1 U901 ( .A1(n4559), .A2(n4560), .A3(n4561), .A4(n4562), .ZN(n4537)
         );
  NAND4_X1 U902 ( .A1(n4539), .A2(n4540), .A3(n4541), .A4(n4542), .ZN(n4538)
         );
  OAI21_X1 U903 ( .B1(n4575), .B2(n4576), .A(n3713), .ZN(n4559) );
  OAI21_X1 U904 ( .B1(n4365), .B2(n4366), .A(n3659), .ZN(n4364) );
  NAND4_X1 U905 ( .A1(n4387), .A2(n4388), .A3(n4389), .A4(n4390), .ZN(n4365)
         );
  NAND4_X1 U906 ( .A1(n4367), .A2(n4368), .A3(n4369), .A4(n4370), .ZN(n4366)
         );
  OAI21_X1 U907 ( .B1(n4403), .B2(n4404), .A(n3713), .ZN(n4387) );
  OAI21_X1 U908 ( .B1(n4193), .B2(n4194), .A(n3659), .ZN(n4192) );
  NAND4_X1 U909 ( .A1(n4215), .A2(n4216), .A3(n4217), .A4(n4218), .ZN(n4193)
         );
  NAND4_X1 U910 ( .A1(n4195), .A2(n4196), .A3(n4197), .A4(n4198), .ZN(n4194)
         );
  OAI21_X1 U911 ( .B1(n4231), .B2(n4232), .A(n3713), .ZN(n4215) );
  OAI21_X1 U912 ( .B1(n4021), .B2(n4022), .A(n3659), .ZN(n4020) );
  NAND4_X1 U913 ( .A1(n4043), .A2(n4044), .A3(n4045), .A4(n4046), .ZN(n4021)
         );
  NAND4_X1 U914 ( .A1(n4023), .A2(n4024), .A3(n4025), .A4(n4026), .ZN(n4022)
         );
  OAI21_X1 U915 ( .B1(n4059), .B2(n4060), .A(n3146), .ZN(n4043) );
  NOR2_X1 U916 ( .A1(n3231), .A2(addr_r[5]), .ZN(n5025) );
  OAI21_X1 U917 ( .B1(n3891), .B2(n3892), .A(n3718), .ZN(n3847) );
  NAND4_X1 U918 ( .A1(n3913), .A2(n3914), .A3(n3915), .A4(n3916), .ZN(n3891)
         );
  NAND4_X1 U919 ( .A1(n3893), .A2(n3894), .A3(n3895), .A4(n3896), .ZN(n3892)
         );
  OAI21_X1 U920 ( .B1(n3929), .B2(n3930), .A(n3713), .ZN(n3913) );
  OAI21_X1 U921 ( .B1(n3716), .B2(n3717), .A(n3718), .ZN(n3655) );
  NAND4_X1 U922 ( .A1(n3739), .A2(n3740), .A3(n3741), .A4(n3742), .ZN(n3716)
         );
  NAND4_X1 U923 ( .A1(n3719), .A2(n3720), .A3(n3721), .A4(n3722), .ZN(n3717)
         );
  OAI21_X1 U924 ( .B1(n3755), .B2(n3756), .A(n3713), .ZN(n3739) );
  AND2_X1 U925 ( .A1(addr_r[3]), .A2(n5015), .ZN(n3698) );
  AND2_X1 U926 ( .A1(n5020), .A2(addr_r[3]), .ZN(n3703) );
  AND2_X1 U927 ( .A1(n5025), .A2(addr_r[3]), .ZN(n3708) );
  AND2_X1 U928 ( .A1(n5030), .A2(addr_r[3]), .ZN(n3713) );
  AND2_X1 U929 ( .A1(addr_r[1]), .A2(n3229), .ZN(n5055) );
  AND2_X1 U930 ( .A1(addr_r[0]), .A2(n5054), .ZN(n3675) );
  AND2_X1 U931 ( .A1(n5052), .A2(addr_r[0]), .ZN(n3670) );
  AND2_X1 U932 ( .A1(addr_r[5]), .A2(addr_r[4]), .ZN(n5015) );
  AND2_X1 U933 ( .A1(addr_r[5]), .A2(n3231), .ZN(n5020) );
  AND2_X1 U934 ( .A1(addr_r[7]), .A2(addr_r[6]), .ZN(n3659) );
  AND2_X1 U935 ( .A1(addr_r[7]), .A2(n3232), .ZN(n3718) );
  INV_X1 U936 ( .A(addr_r[6]), .ZN(n3232) );
  NOR2_X1 U937 ( .A1(n7245), .A2(addr_w[0]), .ZN(n3639) );
  NOR2_X1 U938 ( .A1(addr_w[0]), .A2(addr_w[1]), .ZN(n3634) );
  NOR2_X1 U939 ( .A1(n7116), .A2(addr_w[1]), .ZN(n3631) );
  NOR2_X1 U940 ( .A1(addr_w[2]), .A2(addr_w[3]), .ZN(n3648) );
  NOR2_X1 U941 ( .A1(n7246), .A2(addr_w[3]), .ZN(n3643) );
  NOR2_X1 U942 ( .A1(n7247), .A2(addr_w[2]), .ZN(n3636) );
  NOR2_X1 U943 ( .A1(addr_w[6]), .A2(addr_w[7]), .ZN(n3489) );
  NOR2_X1 U944 ( .A1(n7248), .A2(addr_w[5]), .ZN(n3454) );
  NOR2_X1 U945 ( .A1(addr_w[4]), .A2(addr_w[5]), .ZN(n3399) );
  NOR2_X1 U946 ( .A1(n7250), .A2(addr_w[6]), .ZN(n3398) );
  AND2_X1 U947 ( .A1(addr_w[5]), .A2(n7248), .ZN(n3436) );
  AND2_X1 U948 ( .A1(addr_w[5]), .A2(addr_w[4]), .ZN(n3417) );
  INV_X1 U949 ( .A(addr_w[1]), .ZN(n7245) );
  INV_X1 U950 ( .A(addr_w[2]), .ZN(n7246) );
  INV_X1 U951 ( .A(addr_w[3]), .ZN(n7247) );
  INV_X1 U952 ( .A(addr_w[0]), .ZN(n7116) );
  INV_X1 U953 ( .A(addr_w[6]), .ZN(n7249) );
  INV_X1 U954 ( .A(addr_w[4]), .ZN(n7248) );
  OAI221_X1 U955 ( .B1(n2688), .B2(n3219), .C1(n2680), .C2(n3668), .A(n4921), 
        .ZN(n4920) );
  AOI22_X1 U956 ( .A1(n3201), .A2(n[993]), .B1(n3193), .B2(n[1001]), .ZN(n4921) );
  OAI221_X1 U957 ( .B1(n2112), .B2(n3220), .C1(n2104), .C2(n3668), .A(n4935), 
        .ZN(n4934) );
  AOI22_X1 U958 ( .A1(n3202), .A2(n[1313]), .B1(n3190), .B2(n[1321]), .ZN(
        n4935) );
  OAI221_X1 U959 ( .B1(n1856), .B2(n3223), .C1(n1848), .C2(n3209), .A(n4939), 
        .ZN(n4938) );
  AOI22_X1 U960 ( .A1(n3202), .A2(n[1441]), .B1(n3190), .B2(n[1449]), .ZN(
        n4939) );
  OAI221_X1 U961 ( .B1(n1600), .B2(n3223), .C1(n1592), .C2(n3209), .A(n4943), 
        .ZN(n4942) );
  AOI22_X1 U962 ( .A1(n3208), .A2(n[1569]), .B1(n3198), .B2(n[1577]), .ZN(
        n4943) );
  OAI221_X1 U963 ( .B1(n2240), .B2(n3226), .C1(n2232), .C2(n3217), .A(n4955), 
        .ZN(n4954) );
  AOI22_X1 U964 ( .A1(n3207), .A2(n[1249]), .B1(n3190), .B2(n[1257]), .ZN(
        n4955) );
  OAI221_X1 U965 ( .B1(n1984), .B2(n3225), .C1(n1976), .C2(n3209), .A(n4959), 
        .ZN(n4958) );
  AOI22_X1 U966 ( .A1(n3201), .A2(n[1377]), .B1(n3194), .B2(n[1385]), .ZN(
        n4959) );
  OAI221_X1 U967 ( .B1(n1728), .B2(n3221), .C1(n1720), .C2(n3209), .A(n4963), 
        .ZN(n4962) );
  AOI22_X1 U968 ( .A1(n3204), .A2(n[1505]), .B1(n3194), .B2(n[1513]), .ZN(
        n4963) );
  OAI221_X1 U969 ( .B1(n1088), .B2(n3219), .C1(n1080), .C2(n3213), .A(n4977), 
        .ZN(n4976) );
  AOI22_X1 U970 ( .A1(n3202), .A2(n[1825]), .B1(n3190), .B2(n[1833]), .ZN(
        n4977) );
  OAI221_X1 U971 ( .B1(n832), .B2(n3222), .C1(n824), .C2(n3209), .A(n4981), 
        .ZN(n4980) );
  AOI22_X1 U972 ( .A1(n3200), .A2(n[1953]), .B1(n3196), .B2(n[1961]), .ZN(
        n4981) );
  OAI221_X1 U973 ( .B1(n576), .B2(n3226), .C1(n568), .C2(n3209), .A(n4985), 
        .ZN(n4984) );
  AOI22_X1 U974 ( .A1(n3204), .A2(n[2081]), .B1(n3193), .B2(n[2089]), .ZN(
        n4985) );
  OAI221_X1 U975 ( .B1(n1216), .B2(n3218), .C1(n1208), .C2(n3213), .A(n4997), 
        .ZN(n4996) );
  AOI22_X1 U976 ( .A1(n3201), .A2(n[1761]), .B1(n3191), .B2(n[1769]), .ZN(
        n4997) );
  OAI221_X1 U977 ( .B1(n960), .B2(n3224), .C1(n952), .C2(n3212), .A(n5001), 
        .ZN(n5000) );
  AOI22_X1 U978 ( .A1(n3205), .A2(n[1889]), .B1(n3191), .B2(n[1897]), .ZN(
        n5001) );
  OAI221_X1 U979 ( .B1(n704), .B2(n3667), .C1(n696), .C2(n3210), .A(n5005), 
        .ZN(n5004) );
  AOI22_X1 U980 ( .A1(n3200), .A2(n[2017]), .B1(n3191), .B2(n[2025]), .ZN(
        n5005) );
  OAI221_X1 U981 ( .B1(n320), .B2(n3223), .C1(n312), .C2(n3216), .A(n5021), 
        .ZN(n5019) );
  AOI22_X1 U982 ( .A1(n3670), .A2(n[2337]), .B1(n3191), .B2(n[2345]), .ZN(
        n5021) );
  OAI221_X1 U983 ( .B1(n192), .B2(n3221), .C1(n184), .C2(n3214), .A(n5026), 
        .ZN(n5024) );
  AOI22_X1 U984 ( .A1(n3203), .A2(n[2465]), .B1(n3191), .B2(n[2473]), .ZN(
        n5026) );
  OAI221_X1 U985 ( .B1(n64), .B2(n3667), .C1(n56), .C2(n3214), .A(n5031), .ZN(
        n5029) );
  AOI22_X1 U986 ( .A1(n3206), .A2(n[2593]), .B1(n3191), .B2(n[2601]), .ZN(
        n5031) );
  OAI221_X1 U987 ( .B1(n384), .B2(n3667), .C1(n376), .C2(n3213), .A(n5043), 
        .ZN(n5042) );
  AOI22_X1 U988 ( .A1(n3208), .A2(n[2273]), .B1(n3191), .B2(n[2281]), .ZN(
        n5043) );
  OAI221_X1 U989 ( .B1(n256), .B2(n3667), .C1(n248), .C2(n3212), .A(n5047), 
        .ZN(n5046) );
  AOI22_X1 U990 ( .A1(n3208), .A2(n[2401]), .B1(n3191), .B2(n[2409]), .ZN(
        n5047) );
  OAI221_X1 U991 ( .B1(n128), .B2(n3667), .C1(n120), .C2(n3215), .A(n5051), 
        .ZN(n5050) );
  AOI22_X1 U992 ( .A1(n3201), .A2(n[2529]), .B1(n3191), .B2(n[2537]), .ZN(
        n5051) );
  OAI221_X1 U993 ( .B1(n2687), .B2(n3225), .C1(n2679), .C2(n3210), .A(n4749), 
        .ZN(n4748) );
  AOI22_X1 U994 ( .A1(n3670), .A2(n[994]), .B1(n3192), .B2(n[1002]), .ZN(n4749) );
  OAI221_X1 U995 ( .B1(n2111), .B2(n3226), .C1(n2103), .C2(n3217), .A(n4763), 
        .ZN(n4762) );
  AOI22_X1 U996 ( .A1(n3199), .A2(n[1314]), .B1(n3191), .B2(n[1322]), .ZN(
        n4763) );
  OAI221_X1 U997 ( .B1(n1855), .B2(n3220), .C1(n1847), .C2(n3209), .A(n4767), 
        .ZN(n4766) );
  AOI22_X1 U998 ( .A1(n3201), .A2(n[1442]), .B1(n3198), .B2(n[1450]), .ZN(
        n4767) );
  OAI221_X1 U999 ( .B1(n1599), .B2(n3223), .C1(n1591), .C2(n3217), .A(n4771), 
        .ZN(n4770) );
  AOI22_X1 U1000 ( .A1(n3204), .A2(n[1570]), .B1(n3198), .B2(n[1578]), .ZN(
        n4771) );
  OAI221_X1 U1001 ( .B1(n2239), .B2(n3225), .C1(n2231), .C2(n3668), .A(n4783), 
        .ZN(n4782) );
  AOI22_X1 U1002 ( .A1(n3203), .A2(n[1250]), .B1(n3190), .B2(n[1258]), .ZN(
        n4783) );
  OAI221_X1 U1003 ( .B1(n1983), .B2(n3221), .C1(n1975), .C2(n3209), .A(n4787), 
        .ZN(n4786) );
  AOI22_X1 U1004 ( .A1(n3201), .A2(n[1378]), .B1(n3671), .B2(n[1386]), .ZN(
        n4787) );
  OAI221_X1 U1005 ( .B1(n1727), .B2(n3219), .C1(n1719), .C2(n3212), .A(n4791), 
        .ZN(n4790) );
  AOI22_X1 U1006 ( .A1(n3670), .A2(n[1506]), .B1(n3192), .B2(n[1514]), .ZN(
        n4791) );
  OAI221_X1 U1007 ( .B1(n1087), .B2(n3225), .C1(n1079), .C2(n3211), .A(n4805), 
        .ZN(n4804) );
  AOI22_X1 U1008 ( .A1(n3207), .A2(n[1826]), .B1(n3192), .B2(n[1834]), .ZN(
        n4805) );
  OAI221_X1 U1009 ( .B1(n831), .B2(n3224), .C1(n823), .C2(n3668), .A(n4809), 
        .ZN(n4808) );
  AOI22_X1 U1010 ( .A1(n3203), .A2(n[1954]), .B1(n3192), .B2(n[1962]), .ZN(
        n4809) );
  OAI221_X1 U1011 ( .B1(n575), .B2(n3220), .C1(n567), .C2(n3210), .A(n4813), 
        .ZN(n4812) );
  AOI22_X1 U1012 ( .A1(n3207), .A2(n[2082]), .B1(n3192), .B2(n[2090]), .ZN(
        n4813) );
  OAI221_X1 U1013 ( .B1(n1215), .B2(n3226), .C1(n1207), .C2(n3211), .A(n4825), 
        .ZN(n4824) );
  AOI22_X1 U1014 ( .A1(n3200), .A2(n[1762]), .B1(n3192), .B2(n[1770]), .ZN(
        n4825) );
  OAI221_X1 U1015 ( .B1(n959), .B2(n3224), .C1(n951), .C2(n3213), .A(n4829), 
        .ZN(n4828) );
  AOI22_X1 U1016 ( .A1(n3203), .A2(n[1890]), .B1(n3192), .B2(n[1898]), .ZN(
        n4829) );
  OAI221_X1 U1017 ( .B1(n703), .B2(n3225), .C1(n695), .C2(n3210), .A(n4833), 
        .ZN(n4832) );
  AOI22_X1 U1018 ( .A1(n3201), .A2(n[2018]), .B1(n3192), .B2(n[2026]), .ZN(
        n4833) );
  OAI221_X1 U1019 ( .B1(n319), .B2(n3219), .C1(n311), .C2(n3668), .A(n4847), 
        .ZN(n4846) );
  AOI22_X1 U1020 ( .A1(n3199), .A2(n[2338]), .B1(n3192), .B2(n[2346]), .ZN(
        n4847) );
  OAI221_X1 U1021 ( .B1(n191), .B2(n3226), .C1(n183), .C2(n3217), .A(n4851), 
        .ZN(n4850) );
  AOI22_X1 U1022 ( .A1(n3200), .A2(n[2466]), .B1(n3192), .B2(n[2474]), .ZN(
        n4851) );
  OAI221_X1 U1023 ( .B1(n63), .B2(n3221), .C1(n55), .C2(n3210), .A(n4855), 
        .ZN(n4854) );
  AOI22_X1 U1024 ( .A1(n3208), .A2(n[2594]), .B1(n3192), .B2(n[2602]), .ZN(
        n4855) );
  OAI221_X1 U1025 ( .B1(n383), .B2(n3220), .C1(n375), .C2(n3668), .A(n4867), 
        .ZN(n4866) );
  AOI22_X1 U1026 ( .A1(n3208), .A2(n[2274]), .B1(n3196), .B2(n[2282]), .ZN(
        n4867) );
  OAI221_X1 U1027 ( .B1(n255), .B2(n3226), .C1(n247), .C2(n3668), .A(n4871), 
        .ZN(n4870) );
  AOI22_X1 U1028 ( .A1(n3204), .A2(n[2402]), .B1(n3198), .B2(n[2410]), .ZN(
        n4871) );
  OAI221_X1 U1029 ( .B1(n127), .B2(n3222), .C1(n119), .C2(n3668), .A(n4875), 
        .ZN(n4874) );
  AOI22_X1 U1030 ( .A1(n3670), .A2(n[2530]), .B1(n3196), .B2(n[2538]), .ZN(
        n4875) );
  OAI221_X1 U1031 ( .B1(n1086), .B2(n3226), .C1(n1078), .C2(n3212), .A(n4633), 
        .ZN(n4632) );
  AOI22_X1 U1032 ( .A1(n3670), .A2(n[1827]), .B1(n3195), .B2(n[1835]), .ZN(
        n4633) );
  OAI221_X1 U1033 ( .B1(n830), .B2(n3226), .C1(n822), .C2(n3214), .A(n4637), 
        .ZN(n4636) );
  AOI22_X1 U1034 ( .A1(n3670), .A2(n[1955]), .B1(n3671), .B2(n[1963]), .ZN(
        n4637) );
  OAI221_X1 U1035 ( .B1(n574), .B2(n3219), .C1(n566), .C2(n3668), .A(n4641), 
        .ZN(n4640) );
  AOI22_X1 U1036 ( .A1(n3208), .A2(n[2083]), .B1(n3197), .B2(n[2091]), .ZN(
        n4641) );
  OAI221_X1 U1037 ( .B1(n1214), .B2(n3222), .C1(n1206), .C2(n3214), .A(n4653), 
        .ZN(n4652) );
  AOI22_X1 U1038 ( .A1(n3204), .A2(n[1763]), .B1(n3195), .B2(n[1771]), .ZN(
        n4653) );
  OAI221_X1 U1039 ( .B1(n958), .B2(n3226), .C1(n950), .C2(n3209), .A(n4657), 
        .ZN(n4656) );
  AOI22_X1 U1040 ( .A1(n3206), .A2(n[1891]), .B1(n3194), .B2(n[1899]), .ZN(
        n4657) );
  OAI221_X1 U1041 ( .B1(n702), .B2(n3222), .C1(n694), .C2(n3210), .A(n4661), 
        .ZN(n4660) );
  AOI22_X1 U1042 ( .A1(n3203), .A2(n[2019]), .B1(n3194), .B2(n[2027]), .ZN(
        n4661) );
  OAI221_X1 U1043 ( .B1(n2238), .B2(n3226), .C1(n2230), .C2(n3209), .A(n4611), 
        .ZN(n4610) );
  AOI22_X1 U1044 ( .A1(n3202), .A2(n[1251]), .B1(n3671), .B2(n[1259]), .ZN(
        n4611) );
  OAI221_X1 U1045 ( .B1(n1982), .B2(n3226), .C1(n1974), .C2(n3217), .A(n4615), 
        .ZN(n4614) );
  AOI22_X1 U1046 ( .A1(n3200), .A2(n[1379]), .B1(n3191), .B2(n[1387]), .ZN(
        n4615) );
  OAI221_X1 U1047 ( .B1(n1726), .B2(n3224), .C1(n1718), .C2(n3211), .A(n4619), 
        .ZN(n4618) );
  AOI22_X1 U1048 ( .A1(n3199), .A2(n[1507]), .B1(n3193), .B2(n[1515]), .ZN(
        n4619) );
  OAI221_X1 U1049 ( .B1(n318), .B2(n3218), .C1(n310), .C2(n3209), .A(n4675), 
        .ZN(n4674) );
  AOI22_X1 U1050 ( .A1(n3208), .A2(n[2339]), .B1(n3198), .B2(n[2347]), .ZN(
        n4675) );
  OAI221_X1 U1051 ( .B1(n190), .B2(n3218), .C1(n182), .C2(n3213), .A(n4679), 
        .ZN(n4678) );
  AOI22_X1 U1052 ( .A1(n3201), .A2(n[2467]), .B1(n3191), .B2(n[2475]), .ZN(
        n4679) );
  OAI221_X1 U1053 ( .B1(n62), .B2(n3218), .C1(n54), .C2(n3216), .A(n4683), 
        .ZN(n4682) );
  AOI22_X1 U1054 ( .A1(n3670), .A2(n[2595]), .B1(n3190), .B2(n[2603]), .ZN(
        n4683) );
  OAI221_X1 U1055 ( .B1(n382), .B2(n3218), .C1(n374), .C2(n3213), .A(n4695), 
        .ZN(n4694) );
  AOI22_X1 U1056 ( .A1(n3670), .A2(n[2275]), .B1(n3197), .B2(n[2283]), .ZN(
        n4695) );
  OAI221_X1 U1057 ( .B1(n254), .B2(n3218), .C1(n246), .C2(n3215), .A(n4699), 
        .ZN(n4698) );
  AOI22_X1 U1058 ( .A1(n3670), .A2(n[2403]), .B1(n3194), .B2(n[2411]), .ZN(
        n4699) );
  OAI221_X1 U1059 ( .B1(n126), .B2(n3218), .C1(n118), .C2(n3214), .A(n4703), 
        .ZN(n4702) );
  AOI22_X1 U1060 ( .A1(n3670), .A2(n[2531]), .B1(n3192), .B2(n[2539]), .ZN(
        n4703) );
  OAI221_X1 U1061 ( .B1(n2684), .B2(n3220), .C1(n2676), .C2(n3211), .A(n4233), 
        .ZN(n4232) );
  AOI22_X1 U1062 ( .A1(n3200), .A2(n[997]), .B1(n3194), .B2(n[1005]), .ZN(
        n4233) );
  OAI221_X1 U1063 ( .B1(n2108), .B2(n3220), .C1(n2100), .C2(n3211), .A(n4247), 
        .ZN(n4246) );
  AOI22_X1 U1064 ( .A1(n3200), .A2(n[1317]), .B1(n3194), .B2(n[1325]), .ZN(
        n4247) );
  OAI221_X1 U1065 ( .B1(n1852), .B2(n3220), .C1(n1844), .C2(n3211), .A(n4251), 
        .ZN(n4250) );
  AOI22_X1 U1066 ( .A1(n3200), .A2(n[1445]), .B1(n3194), .B2(n[1453]), .ZN(
        n4251) );
  OAI221_X1 U1067 ( .B1(n1596), .B2(n3220), .C1(n1588), .C2(n3211), .A(n4255), 
        .ZN(n4254) );
  AOI22_X1 U1068 ( .A1(n3200), .A2(n[1573]), .B1(n3194), .B2(n[1581]), .ZN(
        n4255) );
  OAI221_X1 U1069 ( .B1(n2236), .B2(n3220), .C1(n2228), .C2(n3211), .A(n4267), 
        .ZN(n4266) );
  AOI22_X1 U1070 ( .A1(n3200), .A2(n[1253]), .B1(n3194), .B2(n[1261]), .ZN(
        n4267) );
  OAI221_X1 U1071 ( .B1(n1980), .B2(n3220), .C1(n1972), .C2(n3211), .A(n4271), 
        .ZN(n4270) );
  AOI22_X1 U1072 ( .A1(n3200), .A2(n[1381]), .B1(n3194), .B2(n[1389]), .ZN(
        n4271) );
  OAI221_X1 U1073 ( .B1(n1724), .B2(n3220), .C1(n1716), .C2(n3211), .A(n4275), 
        .ZN(n4274) );
  AOI22_X1 U1074 ( .A1(n3200), .A2(n[1509]), .B1(n3194), .B2(n[1517]), .ZN(
        n4275) );
  OAI221_X1 U1075 ( .B1(n1084), .B2(n3219), .C1(n1076), .C2(n3210), .A(n4289), 
        .ZN(n4288) );
  AOI22_X1 U1076 ( .A1(n3199), .A2(n[1829]), .B1(n3193), .B2(n[1837]), .ZN(
        n4289) );
  OAI221_X1 U1077 ( .B1(n828), .B2(n3219), .C1(n820), .C2(n3210), .A(n4293), 
        .ZN(n4292) );
  AOI22_X1 U1078 ( .A1(n3199), .A2(n[1957]), .B1(n3193), .B2(n[1965]), .ZN(
        n4293) );
  OAI221_X1 U1079 ( .B1(n572), .B2(n3219), .C1(n564), .C2(n3210), .A(n4297), 
        .ZN(n4296) );
  AOI22_X1 U1080 ( .A1(n3199), .A2(n[2085]), .B1(n3193), .B2(n[2093]), .ZN(
        n4297) );
  OAI221_X1 U1081 ( .B1(n1212), .B2(n3219), .C1(n1204), .C2(n3210), .A(n4309), 
        .ZN(n4308) );
  AOI22_X1 U1082 ( .A1(n3199), .A2(n[1765]), .B1(n3193), .B2(n[1773]), .ZN(
        n4309) );
  OAI221_X1 U1083 ( .B1(n956), .B2(n3219), .C1(n948), .C2(n3210), .A(n4313), 
        .ZN(n4312) );
  AOI22_X1 U1084 ( .A1(n3199), .A2(n[1893]), .B1(n3193), .B2(n[1901]), .ZN(
        n4313) );
  OAI221_X1 U1085 ( .B1(n700), .B2(n3219), .C1(n692), .C2(n3210), .A(n4317), 
        .ZN(n4316) );
  AOI22_X1 U1086 ( .A1(n3199), .A2(n[2021]), .B1(n3193), .B2(n[2029]), .ZN(
        n4317) );
  OAI221_X1 U1087 ( .B1(n316), .B2(n3219), .C1(n308), .C2(n3210), .A(n4331), 
        .ZN(n4330) );
  AOI22_X1 U1088 ( .A1(n3199), .A2(n[2341]), .B1(n3193), .B2(n[2349]), .ZN(
        n4331) );
  OAI221_X1 U1089 ( .B1(n188), .B2(n3219), .C1(n180), .C2(n3210), .A(n4335), 
        .ZN(n4334) );
  AOI22_X1 U1090 ( .A1(n3199), .A2(n[2469]), .B1(n3193), .B2(n[2477]), .ZN(
        n4335) );
  OAI221_X1 U1091 ( .B1(n60), .B2(n3219), .C1(n52), .C2(n3210), .A(n4339), 
        .ZN(n4338) );
  AOI22_X1 U1092 ( .A1(n3199), .A2(n[2597]), .B1(n3193), .B2(n[2605]), .ZN(
        n4339) );
  OAI221_X1 U1093 ( .B1(n2683), .B2(n3223), .C1(n2675), .C2(n3211), .A(n4061), 
        .ZN(n4060) );
  AOI22_X1 U1094 ( .A1(n3203), .A2(n[998]), .B1(n3197), .B2(n[1006]), .ZN(
        n4061) );
  OAI221_X1 U1095 ( .B1(n2107), .B2(n3223), .C1(n2099), .C2(n3211), .A(n4075), 
        .ZN(n4074) );
  AOI22_X1 U1096 ( .A1(n3203), .A2(n[1318]), .B1(n3197), .B2(n[1326]), .ZN(
        n4075) );
  OAI221_X1 U1097 ( .B1(n1851), .B2(n3223), .C1(n1843), .C2(n3215), .A(n4079), 
        .ZN(n4078) );
  AOI22_X1 U1098 ( .A1(n3203), .A2(n[1446]), .B1(n3197), .B2(n[1454]), .ZN(
        n4079) );
  OAI221_X1 U1099 ( .B1(n1595), .B2(n3223), .C1(n1587), .C2(n3215), .A(n4083), 
        .ZN(n4082) );
  AOI22_X1 U1100 ( .A1(n3203), .A2(n[1574]), .B1(n3197), .B2(n[1582]), .ZN(
        n4083) );
  OAI221_X1 U1101 ( .B1(n2235), .B2(n3222), .C1(n2227), .C2(n3214), .A(n4095), 
        .ZN(n4094) );
  AOI22_X1 U1102 ( .A1(n3202), .A2(n[1254]), .B1(n3196), .B2(n[1262]), .ZN(
        n4095) );
  OAI221_X1 U1103 ( .B1(n1979), .B2(n3222), .C1(n1971), .C2(n3212), .A(n4099), 
        .ZN(n4098) );
  AOI22_X1 U1104 ( .A1(n3202), .A2(n[1382]), .B1(n3196), .B2(n[1390]), .ZN(
        n4099) );
  OAI221_X1 U1105 ( .B1(n1723), .B2(n3222), .C1(n1715), .C2(n3215), .A(n4103), 
        .ZN(n4102) );
  AOI22_X1 U1106 ( .A1(n3202), .A2(n[1510]), .B1(n3196), .B2(n[1518]), .ZN(
        n4103) );
  OAI221_X1 U1107 ( .B1(n1083), .B2(n3222), .C1(n1075), .C2(n3210), .A(n4117), 
        .ZN(n4116) );
  AOI22_X1 U1108 ( .A1(n3202), .A2(n[1830]), .B1(n3196), .B2(n[1838]), .ZN(
        n4117) );
  OAI221_X1 U1109 ( .B1(n827), .B2(n3222), .C1(n819), .C2(n3216), .A(n4121), 
        .ZN(n4120) );
  AOI22_X1 U1110 ( .A1(n3202), .A2(n[1958]), .B1(n3196), .B2(n[1966]), .ZN(
        n4121) );
  OAI221_X1 U1111 ( .B1(n571), .B2(n3222), .C1(n563), .C2(n3213), .A(n4125), 
        .ZN(n4124) );
  AOI22_X1 U1112 ( .A1(n3202), .A2(n[2086]), .B1(n3196), .B2(n[2094]), .ZN(
        n4125) );
  OAI221_X1 U1113 ( .B1(n1211), .B2(n3222), .C1(n1203), .C2(n3211), .A(n4137), 
        .ZN(n4136) );
  AOI22_X1 U1114 ( .A1(n3202), .A2(n[1766]), .B1(n3196), .B2(n[1774]), .ZN(
        n4137) );
  OAI221_X1 U1115 ( .B1(n955), .B2(n3222), .C1(n947), .C2(n3214), .A(n4141), 
        .ZN(n4140) );
  AOI22_X1 U1116 ( .A1(n3202), .A2(n[1894]), .B1(n3196), .B2(n[1902]), .ZN(
        n4141) );
  OAI221_X1 U1117 ( .B1(n699), .B2(n3222), .C1(n691), .C2(n3211), .A(n4145), 
        .ZN(n4144) );
  AOI22_X1 U1118 ( .A1(n3202), .A2(n[2022]), .B1(n3196), .B2(n[2030]), .ZN(
        n4145) );
  OAI221_X1 U1119 ( .B1(n315), .B2(n3221), .C1(n307), .C2(n3210), .A(n4159), 
        .ZN(n4158) );
  AOI22_X1 U1120 ( .A1(n3201), .A2(n[2342]), .B1(n3195), .B2(n[2350]), .ZN(
        n4159) );
  OAI221_X1 U1121 ( .B1(n187), .B2(n3221), .C1(n179), .C2(n3212), .A(n4163), 
        .ZN(n4162) );
  AOI22_X1 U1122 ( .A1(n3201), .A2(n[2470]), .B1(n3195), .B2(n[2478]), .ZN(
        n4163) );
  OAI221_X1 U1123 ( .B1(n59), .B2(n3221), .C1(n51), .C2(n3215), .A(n4167), 
        .ZN(n4166) );
  AOI22_X1 U1124 ( .A1(n3201), .A2(n[2598]), .B1(n3195), .B2(n[2606]), .ZN(
        n4167) );
  OAI221_X1 U1125 ( .B1(n379), .B2(n3221), .C1(n371), .C2(n3217), .A(n4179), 
        .ZN(n4178) );
  AOI22_X1 U1126 ( .A1(n3201), .A2(n[2278]), .B1(n3195), .B2(n[2286]), .ZN(
        n4179) );
  OAI221_X1 U1127 ( .B1(n251), .B2(n3221), .C1(n243), .C2(n3211), .A(n4183), 
        .ZN(n4182) );
  AOI22_X1 U1128 ( .A1(n3201), .A2(n[2406]), .B1(n3195), .B2(n[2414]), .ZN(
        n4183) );
  OAI221_X1 U1129 ( .B1(n123), .B2(n3221), .C1(n115), .C2(n3214), .A(n4187), 
        .ZN(n4186) );
  AOI22_X1 U1130 ( .A1(n3201), .A2(n[2534]), .B1(n3195), .B2(n[2542]), .ZN(
        n4187) );
  OAI221_X1 U1131 ( .B1(n1210), .B2(n3224), .C1(n1202), .C2(n3212), .A(n3965), 
        .ZN(n3964) );
  AOI22_X1 U1132 ( .A1(n3204), .A2(n[1767]), .B1(n3198), .B2(n[1775]), .ZN(
        n3965) );
  OAI221_X1 U1133 ( .B1(n954), .B2(n3224), .C1(n946), .C2(n3212), .A(n3969), 
        .ZN(n3968) );
  AOI22_X1 U1134 ( .A1(n3204), .A2(n[1895]), .B1(n3198), .B2(n[1903]), .ZN(
        n3969) );
  OAI221_X1 U1135 ( .B1(n698), .B2(n3224), .C1(n690), .C2(n3212), .A(n3973), 
        .ZN(n3972) );
  AOI22_X1 U1136 ( .A1(n3204), .A2(n[2023]), .B1(n3198), .B2(n[2031]), .ZN(
        n3973) );
  OAI221_X1 U1137 ( .B1(n314), .B2(n3224), .C1(n306), .C2(n3212), .A(n3987), 
        .ZN(n3986) );
  AOI22_X1 U1138 ( .A1(n3204), .A2(n[2343]), .B1(n3198), .B2(n[2351]), .ZN(
        n3987) );
  OAI221_X1 U1139 ( .B1(n186), .B2(n3224), .C1(n178), .C2(n3212), .A(n3991), 
        .ZN(n3990) );
  AOI22_X1 U1140 ( .A1(n3204), .A2(n[2471]), .B1(n3198), .B2(n[2479]), .ZN(
        n3991) );
  OAI221_X1 U1141 ( .B1(n58), .B2(n3224), .C1(n50), .C2(n3212), .A(n3995), 
        .ZN(n3994) );
  AOI22_X1 U1142 ( .A1(n3204), .A2(n[2599]), .B1(n3198), .B2(n[2607]), .ZN(
        n3995) );
  OAI221_X1 U1143 ( .B1(n378), .B2(n3224), .C1(n370), .C2(n3212), .A(n4007), 
        .ZN(n4006) );
  AOI22_X1 U1144 ( .A1(n3204), .A2(n[2279]), .B1(n3198), .B2(n[2287]), .ZN(
        n4007) );
  OAI221_X1 U1145 ( .B1(n250), .B2(n3224), .C1(n242), .C2(n3212), .A(n4011), 
        .ZN(n4010) );
  AOI22_X1 U1146 ( .A1(n3204), .A2(n[2407]), .B1(n3198), .B2(n[2415]), .ZN(
        n4011) );
  OAI221_X1 U1147 ( .B1(n122), .B2(n3224), .C1(n114), .C2(n3212), .A(n4015), 
        .ZN(n4014) );
  AOI22_X1 U1148 ( .A1(n3204), .A2(n[2535]), .B1(n3198), .B2(n[2543]), .ZN(
        n4015) );
  OAI21_X1 U1149 ( .B1(n4895), .B2(n4896), .A(n3151), .ZN(n4884) );
  OAI221_X1 U1150 ( .B1(n2720), .B2(n3186), .C1(n2712), .C2(n3673), .A(n4898), 
        .ZN(n4895) );
  OAI221_X1 U1151 ( .B1(n2752), .B2(n3223), .C1(n2744), .C2(n3668), .A(n4897), 
        .ZN(n4896) );
  AOI22_X1 U1152 ( .A1(n3166), .A2(n[897]), .B1(n3153), .B2(n[905]), .ZN(n4898) );
  OAI21_X1 U1153 ( .B1(n4915), .B2(n4916), .A(n3147), .ZN(n4904) );
  OAI221_X1 U1154 ( .B1(n2784), .B2(n3188), .C1(n2776), .C2(n3673), .A(n4918), 
        .ZN(n4915) );
  OAI221_X1 U1155 ( .B1(n2816), .B2(n3222), .C1(n2808), .C2(n3668), .A(n4917), 
        .ZN(n4916) );
  AOI22_X1 U1156 ( .A1(n3162), .A2(n[833]), .B1(n3153), .B2(n[841]), .ZN(n4918) );
  OAI21_X1 U1157 ( .B1(n4723), .B2(n4724), .A(n3151), .ZN(n4712) );
  OAI221_X1 U1158 ( .B1(n2719), .B2(n3187), .C1(n2711), .C2(n3673), .A(n4726), 
        .ZN(n4723) );
  OAI221_X1 U1159 ( .B1(n2751), .B2(n3218), .C1(n2743), .C2(n3213), .A(n4725), 
        .ZN(n4724) );
  AOI22_X1 U1160 ( .A1(n3169), .A2(n[898]), .B1(n3157), .B2(n[906]), .ZN(n4726) );
  OAI21_X1 U1161 ( .B1(n4743), .B2(n4744), .A(n3147), .ZN(n4732) );
  OAI221_X1 U1162 ( .B1(n2783), .B2(n3182), .C1(n2775), .C2(n3177), .A(n4746), 
        .ZN(n4743) );
  OAI221_X1 U1163 ( .B1(n2815), .B2(n3219), .C1(n2807), .C2(n3210), .A(n4745), 
        .ZN(n4744) );
  AOI22_X1 U1164 ( .A1(n3165), .A2(n[834]), .B1(n3153), .B2(n[842]), .ZN(n4746) );
  OAI21_X1 U1165 ( .B1(n4207), .B2(n4208), .A(n3684), .ZN(n4196) );
  OAI221_X1 U1166 ( .B1(n2716), .B2(n3186), .C1(n2708), .C2(n3173), .A(n4210), 
        .ZN(n4207) );
  OAI221_X1 U1167 ( .B1(n2748), .B2(n3221), .C1(n2740), .C2(n3212), .A(n4209), 
        .ZN(n4208) );
  AOI22_X1 U1168 ( .A1(n3164), .A2(n[901]), .B1(n3157), .B2(n[909]), .ZN(n4210) );
  OAI21_X1 U1169 ( .B1(n4227), .B2(n4228), .A(n3708), .ZN(n4216) );
  OAI221_X1 U1170 ( .B1(n2780), .B2(n3185), .C1(n2772), .C2(n3174), .A(n4230), 
        .ZN(n4227) );
  OAI221_X1 U1171 ( .B1(n2812), .B2(n3220), .C1(n2804), .C2(n3211), .A(n4229), 
        .ZN(n4228) );
  AOI22_X1 U1172 ( .A1(n3163), .A2(n[837]), .B1(n3155), .B2(n[845]), .ZN(n4230) );
  OAI21_X1 U1173 ( .B1(n4035), .B2(n4036), .A(n3151), .ZN(n4024) );
  OAI221_X1 U1174 ( .B1(n2715), .B2(n3188), .C1(n2707), .C2(n3180), .A(n4038), 
        .ZN(n4035) );
  OAI221_X1 U1175 ( .B1(n2747), .B2(n3223), .C1(n2739), .C2(n3210), .A(n4037), 
        .ZN(n4036) );
  AOI22_X1 U1176 ( .A1(n3166), .A2(n[902]), .B1(n3154), .B2(n[910]), .ZN(n4038) );
  OAI21_X1 U1177 ( .B1(n4055), .B2(n4056), .A(n3147), .ZN(n4044) );
  OAI221_X1 U1178 ( .B1(n2779), .B2(n3188), .C1(n2771), .C2(n3178), .A(n4058), 
        .ZN(n4055) );
  OAI221_X1 U1179 ( .B1(n2811), .B2(n3223), .C1(n2803), .C2(n3211), .A(n4057), 
        .ZN(n4056) );
  AOI22_X1 U1180 ( .A1(n3166), .A2(n[838]), .B1(n3161), .B2(n[846]), .ZN(n4058) );
  OAI221_X1 U1181 ( .B1(n2656), .B2(n3186), .C1(n2648), .C2(n3673), .A(n4922), 
        .ZN(n4919) );
  AOI22_X1 U1182 ( .A1(n3165), .A2(n[961]), .B1(n3153), .B2(n[969]), .ZN(n4922) );
  OAI221_X1 U1183 ( .B1(n2048), .B2(n3186), .C1(n2040), .C2(n3176), .A(n4936), 
        .ZN(n4933) );
  AOI22_X1 U1184 ( .A1(n3167), .A2(n[1281]), .B1(n3153), .B2(n[1289]), .ZN(
        n4936) );
  OAI221_X1 U1185 ( .B1(n1792), .B2(n3188), .C1(n1784), .C2(n3172), .A(n4940), 
        .ZN(n4937) );
  AOI22_X1 U1186 ( .A1(n3171), .A2(n[1409]), .B1(n3158), .B2(n[1417]), .ZN(
        n4940) );
  OAI221_X1 U1187 ( .B1(n1536), .B2(n3189), .C1(n1528), .C2(n3172), .A(n4944), 
        .ZN(n4941) );
  AOI22_X1 U1188 ( .A1(n3165), .A2(n[1537]), .B1(n3155), .B2(n[1545]), .ZN(
        n4944) );
  OAI221_X1 U1189 ( .B1(n2176), .B2(n3189), .C1(n2168), .C2(n3172), .A(n4956), 
        .ZN(n4953) );
  AOI22_X1 U1190 ( .A1(n3168), .A2(n[1217]), .B1(n3154), .B2(n[1225]), .ZN(
        n4956) );
  OAI221_X1 U1191 ( .B1(n1920), .B2(n3185), .C1(n1912), .C2(n3172), .A(n4960), 
        .ZN(n4957) );
  AOI22_X1 U1192 ( .A1(n3162), .A2(n[1345]), .B1(n3154), .B2(n[1353]), .ZN(
        n4960) );
  OAI221_X1 U1193 ( .B1(n1664), .B2(n3186), .C1(n1656), .C2(n3172), .A(n4964), 
        .ZN(n4961) );
  AOI22_X1 U1194 ( .A1(n3164), .A2(n[1473]), .B1(n3155), .B2(n[1481]), .ZN(
        n4964) );
  OAI221_X1 U1195 ( .B1(n1024), .B2(n3187), .C1(n1016), .C2(n3172), .A(n4978), 
        .ZN(n4975) );
  AOI22_X1 U1196 ( .A1(n3167), .A2(n[1793]), .B1(n3158), .B2(n[1801]), .ZN(
        n4978) );
  OAI221_X1 U1197 ( .B1(n768), .B2(n3187), .C1(n760), .C2(n3172), .A(n4982), 
        .ZN(n4979) );
  AOI22_X1 U1198 ( .A1(n3163), .A2(n[1921]), .B1(n3159), .B2(n[1929]), .ZN(
        n4982) );
  OAI221_X1 U1199 ( .B1(n544), .B2(n3187), .C1(n536), .C2(n3172), .A(n4986), 
        .ZN(n4983) );
  AOI22_X1 U1200 ( .A1(n3169), .A2(n[2049]), .B1(n3159), .B2(n[2057]), .ZN(
        n4986) );
  OAI221_X1 U1201 ( .B1(n1152), .B2(n3182), .C1(n1144), .C2(n3173), .A(n4998), 
        .ZN(n4995) );
  AOI22_X1 U1202 ( .A1(n3170), .A2(n[1729]), .B1(n3155), .B2(n[1737]), .ZN(
        n4998) );
  OAI221_X1 U1203 ( .B1(n896), .B2(n3182), .C1(n888), .C2(n3174), .A(n5002), 
        .ZN(n4999) );
  AOI22_X1 U1204 ( .A1(n3675), .A2(n[1857]), .B1(n3161), .B2(n[1865]), .ZN(
        n5002) );
  OAI221_X1 U1205 ( .B1(n640), .B2(n3182), .C1(n632), .C2(n3180), .A(n5006), 
        .ZN(n5003) );
  AOI22_X1 U1206 ( .A1(n3169), .A2(n[1985]), .B1(n3156), .B2(n[1993]), .ZN(
        n5006) );
  OAI221_X1 U1207 ( .B1(n288), .B2(n3182), .C1(n280), .C2(n3173), .A(n5022), 
        .ZN(n5018) );
  AOI22_X1 U1208 ( .A1(n3169), .A2(n[2305]), .B1(n3157), .B2(n[2313]), .ZN(
        n5022) );
  OAI221_X1 U1209 ( .B1(n160), .B2(n3182), .C1(n152), .C2(n3173), .A(n5027), 
        .ZN(n5023) );
  AOI22_X1 U1210 ( .A1(n3167), .A2(n[2433]), .B1(n3154), .B2(n[2441]), .ZN(
        n5027) );
  OAI221_X1 U1211 ( .B1(n32), .B2(n3182), .C1(n24), .C2(n3180), .A(n5032), 
        .ZN(n5028) );
  AOI22_X1 U1212 ( .A1(n3170), .A2(n[2561]), .B1(n3160), .B2(n[2569]), .ZN(
        n5032) );
  OAI221_X1 U1213 ( .B1(n352), .B2(n3182), .C1(n344), .C2(n3177), .A(n5044), 
        .ZN(n5041) );
  AOI22_X1 U1214 ( .A1(n3164), .A2(n[2241]), .B1(n3158), .B2(n[2249]), .ZN(
        n5044) );
  OAI221_X1 U1215 ( .B1(n224), .B2(n3182), .C1(n216), .C2(n3175), .A(n5048), 
        .ZN(n5045) );
  AOI22_X1 U1216 ( .A1(n3166), .A2(n[2369]), .B1(n3155), .B2(n[2377]), .ZN(
        n5048) );
  OAI221_X1 U1217 ( .B1(n96), .B2(n3182), .C1(n88), .C2(n3174), .A(n5053), 
        .ZN(n5049) );
  AOI22_X1 U1218 ( .A1(n3163), .A2(n[2497]), .B1(n3157), .B2(n[2505]), .ZN(
        n5053) );
  OAI221_X1 U1219 ( .B1(n2655), .B2(n3189), .C1(n2647), .C2(n3179), .A(n4750), 
        .ZN(n4747) );
  AOI22_X1 U1220 ( .A1(n3675), .A2(n[962]), .B1(n3153), .B2(n[970]), .ZN(n4750) );
  OAI221_X1 U1221 ( .B1(n2047), .B2(n3182), .C1(n2039), .C2(n3172), .A(n4764), 
        .ZN(n4761) );
  AOI22_X1 U1222 ( .A1(n3165), .A2(n[1282]), .B1(n3676), .B2(n[1290]), .ZN(
        n4764) );
  OAI221_X1 U1223 ( .B1(n1791), .B2(n3183), .C1(n1783), .C2(n3180), .A(n4768), 
        .ZN(n4765) );
  AOI22_X1 U1224 ( .A1(n3171), .A2(n[1410]), .B1(n3676), .B2(n[1418]), .ZN(
        n4768) );
  OAI221_X1 U1225 ( .B1(n1535), .B2(n3184), .C1(n1527), .C2(n3172), .A(n4772), 
        .ZN(n4769) );
  AOI22_X1 U1226 ( .A1(n3675), .A2(n[1538]), .B1(n3156), .B2(n[1546]), .ZN(
        n4772) );
  OAI221_X1 U1227 ( .B1(n2175), .B2(n3185), .C1(n2167), .C2(n3673), .A(n4784), 
        .ZN(n4781) );
  AOI22_X1 U1228 ( .A1(n3166), .A2(n[1218]), .B1(n3676), .B2(n[1226]), .ZN(
        n4784) );
  OAI221_X1 U1229 ( .B1(n1919), .B2(n3183), .C1(n1911), .C2(n3176), .A(n4788), 
        .ZN(n4785) );
  AOI22_X1 U1230 ( .A1(n3171), .A2(n[1346]), .B1(n3160), .B2(n[1354]), .ZN(
        n4788) );
  OAI221_X1 U1231 ( .B1(n1663), .B2(n3672), .C1(n1655), .C2(n3176), .A(n4792), 
        .ZN(n4789) );
  AOI22_X1 U1232 ( .A1(n3675), .A2(n[1474]), .B1(n3159), .B2(n[1482]), .ZN(
        n4792) );
  OAI221_X1 U1233 ( .B1(n1023), .B2(n3183), .C1(n1015), .C2(n3178), .A(n4806), 
        .ZN(n4803) );
  AOI22_X1 U1234 ( .A1(n3171), .A2(n[1794]), .B1(n3676), .B2(n[1802]), .ZN(
        n4806) );
  OAI221_X1 U1235 ( .B1(n767), .B2(n3183), .C1(n759), .C2(n3673), .A(n4810), 
        .ZN(n4807) );
  AOI22_X1 U1236 ( .A1(n3166), .A2(n[1922]), .B1(n3676), .B2(n[1930]), .ZN(
        n4810) );
  OAI221_X1 U1237 ( .B1(n543), .B2(n3183), .C1(n535), .C2(n3173), .A(n4814), 
        .ZN(n4811) );
  AOI22_X1 U1238 ( .A1(n3167), .A2(n[2050]), .B1(n3676), .B2(n[2058]), .ZN(
        n4814) );
  OAI221_X1 U1239 ( .B1(n1151), .B2(n3183), .C1(n1143), .C2(n3173), .A(n4826), 
        .ZN(n4823) );
  AOI22_X1 U1240 ( .A1(n3163), .A2(n[1730]), .B1(n3676), .B2(n[1738]), .ZN(
        n4826) );
  OAI221_X1 U1241 ( .B1(n895), .B2(n3183), .C1(n887), .C2(n3179), .A(n4830), 
        .ZN(n4827) );
  AOI22_X1 U1242 ( .A1(n3168), .A2(n[1858]), .B1(n3676), .B2(n[1866]), .ZN(
        n4830) );
  OAI221_X1 U1243 ( .B1(n639), .B2(n3183), .C1(n631), .C2(n3673), .A(n4834), 
        .ZN(n4831) );
  AOI22_X1 U1244 ( .A1(n3169), .A2(n[1986]), .B1(n3676), .B2(n[1994]), .ZN(
        n4834) );
  OAI221_X1 U1245 ( .B1(n287), .B2(n3183), .C1(n279), .C2(n3673), .A(n4848), 
        .ZN(n4845) );
  AOI22_X1 U1246 ( .A1(n3163), .A2(n[2306]), .B1(n3676), .B2(n[2314]), .ZN(
        n4848) );
  OAI221_X1 U1247 ( .B1(n159), .B2(n3183), .C1(n151), .C2(n3673), .A(n4852), 
        .ZN(n4849) );
  AOI22_X1 U1248 ( .A1(n3165), .A2(n[2434]), .B1(n3676), .B2(n[2442]), .ZN(
        n4852) );
  OAI221_X1 U1249 ( .B1(n31), .B2(n3183), .C1(n23), .C2(n3673), .A(n4856), 
        .ZN(n4853) );
  AOI22_X1 U1250 ( .A1(n3162), .A2(n[2562]), .B1(n3676), .B2(n[2570]), .ZN(
        n4856) );
  OAI221_X1 U1251 ( .B1(n351), .B2(n3187), .C1(n343), .C2(n3673), .A(n4868), 
        .ZN(n4865) );
  AOI22_X1 U1252 ( .A1(n3162), .A2(n[2242]), .B1(n3153), .B2(n[2250]), .ZN(
        n4868) );
  OAI221_X1 U1253 ( .B1(n223), .B2(n3189), .C1(n215), .C2(n3173), .A(n4872), 
        .ZN(n4869) );
  AOI22_X1 U1254 ( .A1(n3675), .A2(n[2370]), .B1(n3153), .B2(n[2378]), .ZN(
        n4872) );
  OAI221_X1 U1255 ( .B1(n95), .B2(n3186), .C1(n87), .C2(n3177), .A(n4876), 
        .ZN(n4873) );
  AOI22_X1 U1256 ( .A1(n3675), .A2(n[2498]), .B1(n3153), .B2(n[2506]), .ZN(
        n4876) );
  OAI221_X1 U1257 ( .B1(n1022), .B2(n3186), .C1(n1014), .C2(n3179), .A(n4634), 
        .ZN(n4631) );
  AOI22_X1 U1258 ( .A1(n3675), .A2(n[1795]), .B1(n3159), .B2(n[1803]), .ZN(
        n4634) );
  OAI221_X1 U1259 ( .B1(n766), .B2(n3184), .C1(n758), .C2(n3174), .A(n4638), 
        .ZN(n4635) );
  AOI22_X1 U1260 ( .A1(n3171), .A2(n[1923]), .B1(n3157), .B2(n[1931]), .ZN(
        n4638) );
  OAI221_X1 U1261 ( .B1(n542), .B2(n3672), .C1(n534), .C2(n3175), .A(n4642), 
        .ZN(n4639) );
  AOI22_X1 U1262 ( .A1(n3162), .A2(n[2051]), .B1(n3156), .B2(n[2059]), .ZN(
        n4642) );
  OAI221_X1 U1263 ( .B1(n1150), .B2(n3672), .C1(n1142), .C2(n3172), .A(n4654), 
        .ZN(n4651) );
  AOI22_X1 U1264 ( .A1(n3166), .A2(n[1731]), .B1(n3157), .B2(n[1739]), .ZN(
        n4654) );
  OAI221_X1 U1265 ( .B1(n894), .B2(n3672), .C1(n886), .C2(n3179), .A(n4658), 
        .ZN(n4655) );
  AOI22_X1 U1266 ( .A1(n3167), .A2(n[1859]), .B1(n3161), .B2(n[1867]), .ZN(
        n4658) );
  OAI221_X1 U1267 ( .B1(n638), .B2(n3672), .C1(n630), .C2(n3179), .A(n4662), 
        .ZN(n4659) );
  AOI22_X1 U1268 ( .A1(n3164), .A2(n[1987]), .B1(n3676), .B2(n[1995]), .ZN(
        n4662) );
  OAI221_X1 U1269 ( .B1(n2174), .B2(n3187), .C1(n2166), .C2(n3172), .A(n4612), 
        .ZN(n4609) );
  AOI22_X1 U1270 ( .A1(n3168), .A2(n[1219]), .B1(n3158), .B2(n[1227]), .ZN(
        n4612) );
  OAI221_X1 U1271 ( .B1(n1918), .B2(n3182), .C1(n1910), .C2(n3673), .A(n4616), 
        .ZN(n4613) );
  AOI22_X1 U1272 ( .A1(n3165), .A2(n[1347]), .B1(n3153), .B2(n[1355]), .ZN(
        n4616) );
  OAI221_X1 U1273 ( .B1(n1662), .B2(n3672), .C1(n1654), .C2(n3180), .A(n4620), 
        .ZN(n4617) );
  AOI22_X1 U1274 ( .A1(n3169), .A2(n[1475]), .B1(n3676), .B2(n[1483]), .ZN(
        n4620) );
  OAI221_X1 U1275 ( .B1(n286), .B2(n3184), .C1(n278), .C2(n3673), .A(n4676), 
        .ZN(n4673) );
  AOI22_X1 U1276 ( .A1(n3165), .A2(n[2307]), .B1(n3676), .B2(n[2315]), .ZN(
        n4676) );
  OAI221_X1 U1277 ( .B1(n158), .B2(n3188), .C1(n150), .C2(n3172), .A(n4680), 
        .ZN(n4677) );
  AOI22_X1 U1278 ( .A1(n3167), .A2(n[2435]), .B1(n3153), .B2(n[2443]), .ZN(
        n4680) );
  OAI221_X1 U1279 ( .B1(n30), .B2(n3189), .C1(n22), .C2(n3176), .A(n4684), 
        .ZN(n4681) );
  AOI22_X1 U1280 ( .A1(n3675), .A2(n[2563]), .B1(n3161), .B2(n[2571]), .ZN(
        n4684) );
  OAI221_X1 U1281 ( .B1(n350), .B2(n3672), .C1(n342), .C2(n3179), .A(n4696), 
        .ZN(n4693) );
  AOI22_X1 U1282 ( .A1(n3675), .A2(n[2243]), .B1(n3160), .B2(n[2251]), .ZN(
        n4696) );
  OAI221_X1 U1283 ( .B1(n222), .B2(n3185), .C1(n214), .C2(n3174), .A(n4700), 
        .ZN(n4697) );
  AOI22_X1 U1284 ( .A1(n3675), .A2(n[2371]), .B1(n3676), .B2(n[2379]), .ZN(
        n4700) );
  OAI221_X1 U1285 ( .B1(n94), .B2(n3183), .C1(n86), .C2(n3673), .A(n4704), 
        .ZN(n4701) );
  AOI22_X1 U1286 ( .A1(n3675), .A2(n[2499]), .B1(n3154), .B2(n[2507]), .ZN(
        n4704) );
  OAI221_X1 U1287 ( .B1(n2652), .B2(n3185), .C1(n2644), .C2(n3174), .A(n4234), 
        .ZN(n4231) );
  AOI22_X1 U1288 ( .A1(n3163), .A2(n[965]), .B1(n3155), .B2(n[973]), .ZN(n4234) );
  OAI221_X1 U1289 ( .B1(n2044), .B2(n3185), .C1(n2036), .C2(n3174), .A(n4248), 
        .ZN(n4245) );
  AOI22_X1 U1290 ( .A1(n3163), .A2(n[1285]), .B1(n3155), .B2(n[1293]), .ZN(
        n4248) );
  OAI221_X1 U1291 ( .B1(n1788), .B2(n3185), .C1(n1780), .C2(n3174), .A(n4252), 
        .ZN(n4249) );
  AOI22_X1 U1292 ( .A1(n3163), .A2(n[1413]), .B1(n3155), .B2(n[1421]), .ZN(
        n4252) );
  OAI221_X1 U1293 ( .B1(n1532), .B2(n3185), .C1(n1524), .C2(n3174), .A(n4256), 
        .ZN(n4253) );
  AOI22_X1 U1294 ( .A1(n3163), .A2(n[1541]), .B1(n3155), .B2(n[1549]), .ZN(
        n4256) );
  OAI221_X1 U1295 ( .B1(n2172), .B2(n3185), .C1(n2164), .C2(n3174), .A(n4268), 
        .ZN(n4265) );
  AOI22_X1 U1296 ( .A1(n3163), .A2(n[1221]), .B1(n3155), .B2(n[1229]), .ZN(
        n4268) );
  OAI221_X1 U1297 ( .B1(n1916), .B2(n3185), .C1(n1908), .C2(n3174), .A(n4272), 
        .ZN(n4269) );
  AOI22_X1 U1298 ( .A1(n3163), .A2(n[1349]), .B1(n3155), .B2(n[1357]), .ZN(
        n4272) );
  OAI221_X1 U1299 ( .B1(n1660), .B2(n3185), .C1(n1652), .C2(n3174), .A(n4276), 
        .ZN(n4273) );
  AOI22_X1 U1300 ( .A1(n3163), .A2(n[1477]), .B1(n3155), .B2(n[1485]), .ZN(
        n4276) );
  OAI221_X1 U1301 ( .B1(n1020), .B2(n3184), .C1(n1012), .C2(n3173), .A(n4290), 
        .ZN(n4287) );
  AOI22_X1 U1302 ( .A1(n3162), .A2(n[1797]), .B1(n3154), .B2(n[1805]), .ZN(
        n4290) );
  OAI221_X1 U1303 ( .B1(n764), .B2(n3184), .C1(n756), .C2(n3173), .A(n4294), 
        .ZN(n4291) );
  AOI22_X1 U1304 ( .A1(n3162), .A2(n[1925]), .B1(n3154), .B2(n[1933]), .ZN(
        n4294) );
  OAI221_X1 U1305 ( .B1(n540), .B2(n3184), .C1(n532), .C2(n3173), .A(n4298), 
        .ZN(n4295) );
  AOI22_X1 U1306 ( .A1(n3162), .A2(n[2053]), .B1(n3154), .B2(n[2061]), .ZN(
        n4298) );
  OAI221_X1 U1307 ( .B1(n1148), .B2(n3184), .C1(n1140), .C2(n3173), .A(n4310), 
        .ZN(n4307) );
  AOI22_X1 U1308 ( .A1(n3162), .A2(n[1733]), .B1(n3154), .B2(n[1741]), .ZN(
        n4310) );
  OAI221_X1 U1309 ( .B1(n892), .B2(n3184), .C1(n884), .C2(n3173), .A(n4314), 
        .ZN(n4311) );
  AOI22_X1 U1310 ( .A1(n3162), .A2(n[1861]), .B1(n3154), .B2(n[1869]), .ZN(
        n4314) );
  OAI221_X1 U1311 ( .B1(n636), .B2(n3184), .C1(n628), .C2(n3173), .A(n4318), 
        .ZN(n4315) );
  AOI22_X1 U1312 ( .A1(n3162), .A2(n[1989]), .B1(n3154), .B2(n[1997]), .ZN(
        n4318) );
  OAI221_X1 U1313 ( .B1(n284), .B2(n3184), .C1(n276), .C2(n3173), .A(n4332), 
        .ZN(n4329) );
  AOI22_X1 U1314 ( .A1(n3162), .A2(n[2309]), .B1(n3154), .B2(n[2317]), .ZN(
        n4332) );
  OAI221_X1 U1315 ( .B1(n156), .B2(n3184), .C1(n148), .C2(n3173), .A(n4336), 
        .ZN(n4333) );
  AOI22_X1 U1316 ( .A1(n3162), .A2(n[2437]), .B1(n3154), .B2(n[2445]), .ZN(
        n4336) );
  OAI221_X1 U1317 ( .B1(n28), .B2(n3184), .C1(n20), .C2(n3173), .A(n4340), 
        .ZN(n4337) );
  AOI22_X1 U1318 ( .A1(n3162), .A2(n[2565]), .B1(n3154), .B2(n[2573]), .ZN(
        n4340) );
  OAI221_X1 U1319 ( .B1(n2651), .B2(n3188), .C1(n2643), .C2(n3178), .A(n4062), 
        .ZN(n4059) );
  AOI22_X1 U1320 ( .A1(n3166), .A2(n[966]), .B1(n3159), .B2(n[974]), .ZN(n4062) );
  OAI221_X1 U1321 ( .B1(n2043), .B2(n3188), .C1(n2035), .C2(n3176), .A(n4076), 
        .ZN(n4073) );
  AOI22_X1 U1322 ( .A1(n3166), .A2(n[1286]), .B1(n3159), .B2(n[1294]), .ZN(
        n4076) );
  OAI221_X1 U1323 ( .B1(n1787), .B2(n3188), .C1(n1779), .C2(n3173), .A(n4080), 
        .ZN(n4077) );
  AOI22_X1 U1324 ( .A1(n3166), .A2(n[1414]), .B1(n3156), .B2(n[1422]), .ZN(
        n4080) );
  OAI221_X1 U1325 ( .B1(n1531), .B2(n3188), .C1(n1523), .C2(n3177), .A(n4084), 
        .ZN(n4081) );
  AOI22_X1 U1326 ( .A1(n3166), .A2(n[1542]), .B1(n3158), .B2(n[1550]), .ZN(
        n4084) );
  OAI221_X1 U1327 ( .B1(n2171), .B2(n3187), .C1(n2163), .C2(n3177), .A(n4096), 
        .ZN(n4093) );
  AOI22_X1 U1328 ( .A1(n3165), .A2(n[1222]), .B1(n3155), .B2(n[1230]), .ZN(
        n4096) );
  OAI221_X1 U1329 ( .B1(n1915), .B2(n3187), .C1(n1907), .C2(n3175), .A(n4100), 
        .ZN(n4097) );
  AOI22_X1 U1330 ( .A1(n3165), .A2(n[1350]), .B1(n3155), .B2(n[1358]), .ZN(
        n4100) );
  OAI221_X1 U1331 ( .B1(n1659), .B2(n3187), .C1(n1651), .C2(n3174), .A(n4104), 
        .ZN(n4101) );
  AOI22_X1 U1332 ( .A1(n3165), .A2(n[1478]), .B1(n3161), .B2(n[1486]), .ZN(
        n4104) );
  OAI221_X1 U1333 ( .B1(n1019), .B2(n3187), .C1(n1011), .C2(n3178), .A(n4118), 
        .ZN(n4115) );
  AOI22_X1 U1334 ( .A1(n3165), .A2(n[1798]), .B1(n3158), .B2(n[1806]), .ZN(
        n4118) );
  OAI221_X1 U1335 ( .B1(n763), .B2(n3187), .C1(n755), .C2(n3179), .A(n4122), 
        .ZN(n4119) );
  AOI22_X1 U1336 ( .A1(n3165), .A2(n[1926]), .B1(n3157), .B2(n[1934]), .ZN(
        n4122) );
  OAI221_X1 U1337 ( .B1(n539), .B2(n3187), .C1(n531), .C2(n3176), .A(n4126), 
        .ZN(n4123) );
  AOI22_X1 U1338 ( .A1(n3165), .A2(n[2054]), .B1(n3157), .B2(n[2062]), .ZN(
        n4126) );
  OAI221_X1 U1339 ( .B1(n1147), .B2(n3187), .C1(n1139), .C2(n3173), .A(n4138), 
        .ZN(n4135) );
  AOI22_X1 U1340 ( .A1(n3165), .A2(n[1734]), .B1(n3154), .B2(n[1742]), .ZN(
        n4138) );
  OAI221_X1 U1341 ( .B1(n891), .B2(n3187), .C1(n883), .C2(n3175), .A(n4142), 
        .ZN(n4139) );
  AOI22_X1 U1342 ( .A1(n3165), .A2(n[1862]), .B1(n3160), .B2(n[1870]), .ZN(
        n4142) );
  OAI221_X1 U1343 ( .B1(n635), .B2(n3187), .C1(n627), .C2(n3175), .A(n4146), 
        .ZN(n4143) );
  AOI22_X1 U1344 ( .A1(n3165), .A2(n[1990]), .B1(n3157), .B2(n[1998]), .ZN(
        n4146) );
  OAI221_X1 U1345 ( .B1(n283), .B2(n3186), .C1(n275), .C2(n3177), .A(n4160), 
        .ZN(n4157) );
  AOI22_X1 U1346 ( .A1(n3164), .A2(n[2310]), .B1(n3156), .B2(n[2318]), .ZN(
        n4160) );
  OAI221_X1 U1347 ( .B1(n155), .B2(n3186), .C1(n147), .C2(n3174), .A(n4164), 
        .ZN(n4161) );
  AOI22_X1 U1348 ( .A1(n3164), .A2(n[2438]), .B1(n3153), .B2(n[2446]), .ZN(
        n4164) );
  OAI221_X1 U1349 ( .B1(n27), .B2(n3186), .C1(n19), .C2(n3179), .A(n4168), 
        .ZN(n4165) );
  AOI22_X1 U1350 ( .A1(n3164), .A2(n[2566]), .B1(n3157), .B2(n[2574]), .ZN(
        n4168) );
  OAI221_X1 U1351 ( .B1(n347), .B2(n3186), .C1(n339), .C2(n3176), .A(n4180), 
        .ZN(n4177) );
  AOI22_X1 U1352 ( .A1(n3164), .A2(n[2246]), .B1(n3154), .B2(n[2254]), .ZN(
        n4180) );
  OAI221_X1 U1353 ( .B1(n219), .B2(n3186), .C1(n211), .C2(n3180), .A(n4184), 
        .ZN(n4181) );
  AOI22_X1 U1354 ( .A1(n3164), .A2(n[2374]), .B1(n3154), .B2(n[2382]), .ZN(
        n4184) );
  OAI221_X1 U1355 ( .B1(n91), .B2(n3186), .C1(n83), .C2(n3174), .A(n4188), 
        .ZN(n4185) );
  AOI22_X1 U1356 ( .A1(n3164), .A2(n[2502]), .B1(n3161), .B2(n[2510]), .ZN(
        n4188) );
  OAI221_X1 U1357 ( .B1(n1146), .B2(n3189), .C1(n1138), .C2(n3175), .A(n3966), 
        .ZN(n3963) );
  AOI22_X1 U1358 ( .A1(n3167), .A2(n[1735]), .B1(n3156), .B2(n[1743]), .ZN(
        n3966) );
  OAI221_X1 U1359 ( .B1(n890), .B2(n3189), .C1(n882), .C2(n3175), .A(n3970), 
        .ZN(n3967) );
  AOI22_X1 U1360 ( .A1(n3167), .A2(n[1863]), .B1(n3156), .B2(n[1871]), .ZN(
        n3970) );
  OAI221_X1 U1361 ( .B1(n634), .B2(n3189), .C1(n626), .C2(n3175), .A(n3974), 
        .ZN(n3971) );
  AOI22_X1 U1362 ( .A1(n3167), .A2(n[1991]), .B1(n3156), .B2(n[1999]), .ZN(
        n3974) );
  OAI221_X1 U1363 ( .B1(n282), .B2(n3189), .C1(n274), .C2(n3175), .A(n3988), 
        .ZN(n3985) );
  AOI22_X1 U1364 ( .A1(n3167), .A2(n[2311]), .B1(n3156), .B2(n[2319]), .ZN(
        n3988) );
  OAI221_X1 U1365 ( .B1(n154), .B2(n3189), .C1(n146), .C2(n3175), .A(n3992), 
        .ZN(n3989) );
  AOI22_X1 U1366 ( .A1(n3167), .A2(n[2439]), .B1(n3156), .B2(n[2447]), .ZN(
        n3992) );
  OAI221_X1 U1367 ( .B1(n26), .B2(n3189), .C1(n18), .C2(n3175), .A(n3996), 
        .ZN(n3993) );
  AOI22_X1 U1368 ( .A1(n3167), .A2(n[2567]), .B1(n3156), .B2(n[2575]), .ZN(
        n3996) );
  OAI221_X1 U1369 ( .B1(n346), .B2(n3189), .C1(n338), .C2(n3175), .A(n4008), 
        .ZN(n4005) );
  AOI22_X1 U1370 ( .A1(n3167), .A2(n[2247]), .B1(n3156), .B2(n[2255]), .ZN(
        n4008) );
  OAI221_X1 U1371 ( .B1(n218), .B2(n3189), .C1(n210), .C2(n3175), .A(n4012), 
        .ZN(n4009) );
  AOI22_X1 U1372 ( .A1(n3167), .A2(n[2375]), .B1(n3156), .B2(n[2383]), .ZN(
        n4012) );
  OAI221_X1 U1373 ( .B1(n90), .B2(n3189), .C1(n82), .C2(n3175), .A(n4016), 
        .ZN(n4013) );
  AOI22_X1 U1374 ( .A1(n3167), .A2(n[2503]), .B1(n3156), .B2(n[2511]), .ZN(
        n4016) );
  AOI22_X1 U1375 ( .A1(n3203), .A2(n[673]), .B1(n3671), .B2(n[681]), .ZN(n4889) );
  AOI22_X1 U1376 ( .A1(n3203), .A2(n[801]), .B1(n3195), .B2(n[809]), .ZN(n4893) );
  AOI22_X1 U1377 ( .A1(n3208), .A2(n[929]), .B1(n3197), .B2(n[937]), .ZN(n4897) );
  AOI22_X1 U1378 ( .A1(n3202), .A2(n[1057]), .B1(n3197), .B2(n[1065]), .ZN(
        n4901) );
  AOI22_X1 U1379 ( .A1(n3200), .A2(n[609]), .B1(n3196), .B2(n[617]), .ZN(n4909) );
  AOI22_X1 U1380 ( .A1(n3199), .A2(n[737]), .B1(n3193), .B2(n[745]), .ZN(n4913) );
  AOI22_X1 U1381 ( .A1(n3206), .A2(n[865]), .B1(n3198), .B2(n[873]), .ZN(n4917) );
  AOI22_X1 U1382 ( .A1(n3670), .A2(n[1185]), .B1(n3190), .B2(n[1193]), .ZN(
        n4931) );
  AOI22_X1 U1383 ( .A1(n3199), .A2(n[1121]), .B1(n3190), .B2(n[1129]), .ZN(
        n4951) );
  AOI22_X1 U1384 ( .A1(n3206), .A2(n[1697]), .B1(n3190), .B2(n[1705]), .ZN(
        n4973) );
  AOI22_X1 U1385 ( .A1(n3208), .A2(n[1633]), .B1(n3191), .B2(n[1641]), .ZN(
        n4993) );
  AOI22_X1 U1386 ( .A1(n3199), .A2(n[2209]), .B1(n3191), .B2(n[2217]), .ZN(
        n5016) );
  AOI22_X1 U1387 ( .A1(n3202), .A2(n[2145]), .B1(n3191), .B2(n[2153]), .ZN(
        n5039) );
  AOI22_X1 U1388 ( .A1(n3670), .A2(n[674]), .B1(n3671), .B2(n[682]), .ZN(n4717) );
  AOI22_X1 U1389 ( .A1(n3200), .A2(n[802]), .B1(n3671), .B2(n[810]), .ZN(n4721) );
  AOI22_X1 U1390 ( .A1(n3207), .A2(n[930]), .B1(n3194), .B2(n[938]), .ZN(n4725) );
  AOI22_X1 U1391 ( .A1(n3206), .A2(n[1058]), .B1(n3193), .B2(n[1066]), .ZN(
        n4729) );
  AOI22_X1 U1392 ( .A1(n3207), .A2(n[610]), .B1(n3191), .B2(n[618]), .ZN(n4737) );
  AOI22_X1 U1393 ( .A1(n3202), .A2(n[738]), .B1(n3192), .B2(n[746]), .ZN(n4741) );
  AOI22_X1 U1394 ( .A1(n3208), .A2(n[866]), .B1(n3191), .B2(n[874]), .ZN(n4745) );
  AOI22_X1 U1395 ( .A1(n3205), .A2(n[1186]), .B1(n3192), .B2(n[1194]), .ZN(
        n4759) );
  AOI22_X1 U1396 ( .A1(n3206), .A2(n[1122]), .B1(n3192), .B2(n[1130]), .ZN(
        n4779) );
  AOI22_X1 U1397 ( .A1(n3208), .A2(n[1698]), .B1(n3192), .B2(n[1706]), .ZN(
        n4801) );
  AOI22_X1 U1398 ( .A1(n3206), .A2(n[1634]), .B1(n3192), .B2(n[1642]), .ZN(
        n4821) );
  AOI22_X1 U1399 ( .A1(n3202), .A2(n[2210]), .B1(n3192), .B2(n[2218]), .ZN(
        n4843) );
  AOI22_X1 U1400 ( .A1(n3204), .A2(n[2146]), .B1(n3195), .B2(n[2154]), .ZN(
        n4863) );
  AOI22_X1 U1401 ( .A1(n3670), .A2(n[1699]), .B1(n3194), .B2(n[1707]), .ZN(
        n4629) );
  AOI22_X1 U1402 ( .A1(n3207), .A2(n[1635]), .B1(n3196), .B2(n[1643]), .ZN(
        n4649) );
  AOI22_X1 U1403 ( .A1(n3670), .A2(n[1123]), .B1(n3190), .B2(n[1131]), .ZN(
        n4607) );
  AOI22_X1 U1404 ( .A1(n3200), .A2(n[2211]), .B1(n3196), .B2(n[2219]), .ZN(
        n4671) );
  AOI22_X1 U1405 ( .A1(n3199), .A2(n[2147]), .B1(n3191), .B2(n[2155]), .ZN(
        n4691) );
  AOI22_X1 U1406 ( .A1(n3201), .A2(n[677]), .B1(n3195), .B2(n[685]), .ZN(n4201) );
  AOI22_X1 U1407 ( .A1(n3201), .A2(n[805]), .B1(n3195), .B2(n[813]), .ZN(n4205) );
  AOI22_X1 U1408 ( .A1(n3201), .A2(n[933]), .B1(n3195), .B2(n[941]), .ZN(n4209) );
  AOI22_X1 U1409 ( .A1(n3201), .A2(n[1061]), .B1(n3195), .B2(n[1069]), .ZN(
        n4213) );
  AOI22_X1 U1410 ( .A1(n3200), .A2(n[613]), .B1(n3194), .B2(n[621]), .ZN(n4221) );
  AOI22_X1 U1411 ( .A1(n3200), .A2(n[741]), .B1(n3194), .B2(n[749]), .ZN(n4225) );
  AOI22_X1 U1412 ( .A1(n3200), .A2(n[869]), .B1(n3194), .B2(n[877]), .ZN(n4229) );
  AOI22_X1 U1413 ( .A1(n3200), .A2(n[1189]), .B1(n3194), .B2(n[1197]), .ZN(
        n4243) );
  AOI22_X1 U1414 ( .A1(n3200), .A2(n[1125]), .B1(n3194), .B2(n[1133]), .ZN(
        n4263) );
  AOI22_X1 U1415 ( .A1(n3199), .A2(n[1701]), .B1(n3193), .B2(n[1709]), .ZN(
        n4285) );
  AOI22_X1 U1416 ( .A1(n3199), .A2(n[1637]), .B1(n3193), .B2(n[1645]), .ZN(
        n4305) );
  AOI22_X1 U1417 ( .A1(n3199), .A2(n[2213]), .B1(n3193), .B2(n[2221]), .ZN(
        n4327) );
  AOI22_X1 U1418 ( .A1(n3203), .A2(n[678]), .B1(n3197), .B2(n[686]), .ZN(n4029) );
  AOI22_X1 U1419 ( .A1(n3203), .A2(n[806]), .B1(n3197), .B2(n[814]), .ZN(n4033) );
  AOI22_X1 U1420 ( .A1(n3203), .A2(n[934]), .B1(n3197), .B2(n[942]), .ZN(n4037) );
  AOI22_X1 U1421 ( .A1(n3203), .A2(n[1062]), .B1(n3197), .B2(n[1070]), .ZN(
        n4041) );
  AOI22_X1 U1422 ( .A1(n3203), .A2(n[614]), .B1(n3197), .B2(n[622]), .ZN(n4049) );
  AOI22_X1 U1423 ( .A1(n3203), .A2(n[742]), .B1(n3197), .B2(n[750]), .ZN(n4053) );
  AOI22_X1 U1424 ( .A1(n3203), .A2(n[870]), .B1(n3197), .B2(n[878]), .ZN(n4057) );
  AOI22_X1 U1425 ( .A1(n3203), .A2(n[1190]), .B1(n3197), .B2(n[1198]), .ZN(
        n4071) );
  AOI22_X1 U1426 ( .A1(n3202), .A2(n[1126]), .B1(n3196), .B2(n[1134]), .ZN(
        n4091) );
  AOI22_X1 U1427 ( .A1(n3202), .A2(n[1702]), .B1(n3196), .B2(n[1710]), .ZN(
        n4113) );
  AOI22_X1 U1428 ( .A1(n3202), .A2(n[1638]), .B1(n3196), .B2(n[1646]), .ZN(
        n4133) );
  AOI22_X1 U1429 ( .A1(n3201), .A2(n[2214]), .B1(n3195), .B2(n[2222]), .ZN(
        n4155) );
  AOI22_X1 U1430 ( .A1(n3201), .A2(n[2150]), .B1(n3195), .B2(n[2158]), .ZN(
        n4175) );
  AOI22_X1 U1431 ( .A1(n3204), .A2(n[1639]), .B1(n3198), .B2(n[1647]), .ZN(
        n3961) );
  AOI22_X1 U1432 ( .A1(n3204), .A2(n[2215]), .B1(n3198), .B2(n[2223]), .ZN(
        n3983) );
  AOI22_X1 U1433 ( .A1(n3204), .A2(n[2151]), .B1(n3198), .B2(n[2159]), .ZN(
        n4003) );
  OAI221_X1 U1434 ( .B1(n2873), .B2(n3226), .C1(n2865), .C2(n3217), .A(n3680), 
        .ZN(n3678) );
  AOI22_X1 U1435 ( .A1(n3208), .A2(n[808]), .B1(n3196), .B2(n[816]), .ZN(n3680) );
  OAI221_X1 U1436 ( .B1(n2745), .B2(n3226), .C1(n2737), .C2(n3217), .A(n3685), 
        .ZN(n3683) );
  AOI22_X1 U1437 ( .A1(n3208), .A2(n[936]), .B1(n3190), .B2(n[944]), .ZN(n3685) );
  OAI221_X1 U1438 ( .B1(n2617), .B2(n3226), .C1(n2609), .C2(n3217), .A(n3690), 
        .ZN(n3688) );
  AOI22_X1 U1439 ( .A1(n3208), .A2(n[1064]), .B1(n3193), .B2(n[1072]), .ZN(
        n3690) );
  OAI221_X1 U1440 ( .B1(n2686), .B2(n3226), .C1(n2678), .C2(n3668), .A(n4577), 
        .ZN(n4576) );
  AOI22_X1 U1441 ( .A1(n3205), .A2(n[995]), .B1(n3198), .B2(n[1003]), .ZN(
        n4577) );
  OAI221_X1 U1442 ( .B1(n2110), .B2(n3226), .C1(n2102), .C2(n3217), .A(n4591), 
        .ZN(n4590) );
  AOI22_X1 U1443 ( .A1(n3205), .A2(n[1315]), .B1(n3195), .B2(n[1323]), .ZN(
        n4591) );
  OAI221_X1 U1444 ( .B1(n1854), .B2(n3220), .C1(n1846), .C2(n3217), .A(n4595), 
        .ZN(n4594) );
  AOI22_X1 U1445 ( .A1(n3205), .A2(n[1443]), .B1(n3197), .B2(n[1451]), .ZN(
        n4595) );
  OAI221_X1 U1446 ( .B1(n1598), .B2(n3221), .C1(n1590), .C2(n3212), .A(n4599), 
        .ZN(n4598) );
  AOI22_X1 U1447 ( .A1(n3205), .A2(n[1571]), .B1(n3197), .B2(n[1579]), .ZN(
        n4599) );
  OAI221_X1 U1448 ( .B1(n2685), .B2(n3223), .C1(n2677), .C2(n3214), .A(n4405), 
        .ZN(n4404) );
  AOI22_X1 U1449 ( .A1(n3202), .A2(n[996]), .B1(n3191), .B2(n[1004]), .ZN(
        n4405) );
  OAI221_X1 U1450 ( .B1(n2109), .B2(n3667), .C1(n2101), .C2(n3215), .A(n4419), 
        .ZN(n4418) );
  AOI22_X1 U1451 ( .A1(n3670), .A2(n[1316]), .B1(n3193), .B2(n[1324]), .ZN(
        n4419) );
  OAI221_X1 U1452 ( .B1(n1853), .B2(n3223), .C1(n1845), .C2(n3216), .A(n4423), 
        .ZN(n4422) );
  AOI22_X1 U1453 ( .A1(n3202), .A2(n[1444]), .B1(n3198), .B2(n[1452]), .ZN(
        n4423) );
  OAI221_X1 U1454 ( .B1(n1597), .B2(n3221), .C1(n1589), .C2(n3215), .A(n4427), 
        .ZN(n4426) );
  AOI22_X1 U1455 ( .A1(n3200), .A2(n[1572]), .B1(n3193), .B2(n[1580]), .ZN(
        n4427) );
  OAI221_X1 U1456 ( .B1(n2237), .B2(n3221), .C1(n2229), .C2(n3212), .A(n4439), 
        .ZN(n4438) );
  AOI22_X1 U1457 ( .A1(n3205), .A2(n[1252]), .B1(n3194), .B2(n[1260]), .ZN(
        n4439) );
  OAI221_X1 U1458 ( .B1(n1981), .B2(n3224), .C1(n1973), .C2(n3216), .A(n4443), 
        .ZN(n4442) );
  AOI22_X1 U1459 ( .A1(n3205), .A2(n[1380]), .B1(n3197), .B2(n[1388]), .ZN(
        n4443) );
  OAI221_X1 U1460 ( .B1(n1725), .B2(n3219), .C1(n1717), .C2(n3216), .A(n4447), 
        .ZN(n4446) );
  AOI22_X1 U1461 ( .A1(n3201), .A2(n[1508]), .B1(n3196), .B2(n[1516]), .ZN(
        n4447) );
  OAI221_X1 U1462 ( .B1(n1085), .B2(n3218), .C1(n1077), .C2(n3214), .A(n4461), 
        .ZN(n4460) );
  AOI22_X1 U1463 ( .A1(n3199), .A2(n[1828]), .B1(n3190), .B2(n[1836]), .ZN(
        n4461) );
  OAI221_X1 U1464 ( .B1(n829), .B2(n3220), .C1(n821), .C2(n3210), .A(n4465), 
        .ZN(n4464) );
  AOI22_X1 U1465 ( .A1(n3203), .A2(n[1956]), .B1(n3193), .B2(n[1964]), .ZN(
        n4465) );
  OAI221_X1 U1466 ( .B1(n573), .B2(n3222), .C1(n565), .C2(n3217), .A(n4469), 
        .ZN(n4468) );
  AOI22_X1 U1467 ( .A1(n3204), .A2(n[2084]), .B1(n3671), .B2(n[2092]), .ZN(
        n4469) );
  OAI221_X1 U1468 ( .B1(n1213), .B2(n3219), .C1(n1205), .C2(n3212), .A(n4481), 
        .ZN(n4480) );
  AOI22_X1 U1469 ( .A1(n3208), .A2(n[1764]), .B1(n3195), .B2(n[1772]), .ZN(
        n4481) );
  OAI221_X1 U1470 ( .B1(n957), .B2(n3222), .C1(n949), .C2(n3211), .A(n4485), 
        .ZN(n4484) );
  AOI22_X1 U1471 ( .A1(n3208), .A2(n[1892]), .B1(n3671), .B2(n[1900]), .ZN(
        n4485) );
  OAI221_X1 U1472 ( .B1(n701), .B2(n3223), .C1(n693), .C2(n3216), .A(n4489), 
        .ZN(n4488) );
  AOI22_X1 U1473 ( .A1(n3207), .A2(n[2020]), .B1(n3198), .B2(n[2028]), .ZN(
        n4489) );
  OAI221_X1 U1474 ( .B1(n317), .B2(n3221), .C1(n309), .C2(n3216), .A(n4503), 
        .ZN(n4502) );
  AOI22_X1 U1475 ( .A1(n3208), .A2(n[2340]), .B1(n3190), .B2(n[2348]), .ZN(
        n4503) );
  OAI221_X1 U1476 ( .B1(n189), .B2(n3222), .C1(n181), .C2(n3210), .A(n4507), 
        .ZN(n4506) );
  AOI22_X1 U1477 ( .A1(n3208), .A2(n[2468]), .B1(n3197), .B2(n[2476]), .ZN(
        n4507) );
  OAI221_X1 U1478 ( .B1(n61), .B2(n3226), .C1(n53), .C2(n3211), .A(n4511), 
        .ZN(n4510) );
  AOI22_X1 U1479 ( .A1(n3208), .A2(n[2596]), .B1(n3197), .B2(n[2604]), .ZN(
        n4511) );
  OAI221_X1 U1480 ( .B1(n381), .B2(n3218), .C1(n373), .C2(n3210), .A(n4523), 
        .ZN(n4522) );
  AOI22_X1 U1481 ( .A1(n3208), .A2(n[2276]), .B1(n3197), .B2(n[2284]), .ZN(
        n4523) );
  OAI221_X1 U1482 ( .B1(n253), .B2(n3218), .C1(n245), .C2(n3217), .A(n4527), 
        .ZN(n4526) );
  AOI22_X1 U1483 ( .A1(n3204), .A2(n[2404]), .B1(n3195), .B2(n[2412]), .ZN(
        n4527) );
  OAI221_X1 U1484 ( .B1(n125), .B2(n3667), .C1(n117), .C2(n3217), .A(n4531), 
        .ZN(n4530) );
  AOI22_X1 U1485 ( .A1(n3204), .A2(n[2532]), .B1(n3194), .B2(n[2540]), .ZN(
        n4531) );
  OAI221_X1 U1486 ( .B1(n380), .B2(n3220), .C1(n372), .C2(n3215), .A(n4351), 
        .ZN(n4350) );
  AOI22_X1 U1487 ( .A1(n3201), .A2(n[2277]), .B1(n3197), .B2(n[2285]), .ZN(
        n4351) );
  OAI221_X1 U1488 ( .B1(n252), .B2(n3224), .C1(n244), .C2(n3209), .A(n4355), 
        .ZN(n4354) );
  AOI22_X1 U1489 ( .A1(n3200), .A2(n[2405]), .B1(n3190), .B2(n[2413]), .ZN(
        n4355) );
  OAI221_X1 U1490 ( .B1(n124), .B2(n3667), .C1(n116), .C2(n3212), .A(n4359), 
        .ZN(n4358) );
  AOI22_X1 U1491 ( .A1(n3207), .A2(n[2533]), .B1(n3194), .B2(n[2541]), .ZN(
        n4359) );
  OAI221_X1 U1492 ( .B1(n1722), .B2(n3220), .C1(n1714), .C2(n3213), .A(n3931), 
        .ZN(n3930) );
  AOI22_X1 U1493 ( .A1(n3203), .A2(n[1511]), .B1(n3191), .B2(n[1519]), .ZN(
        n3931) );
  OAI221_X1 U1494 ( .B1(n1082), .B2(n3220), .C1(n1074), .C2(n3213), .A(n3945), 
        .ZN(n3944) );
  AOI22_X1 U1495 ( .A1(n3200), .A2(n[1831]), .B1(n3191), .B2(n[1839]), .ZN(
        n3945) );
  OAI221_X1 U1496 ( .B1(n826), .B2(n3220), .C1(n818), .C2(n3213), .A(n3949), 
        .ZN(n3948) );
  AOI22_X1 U1497 ( .A1(n3206), .A2(n[1959]), .B1(n3195), .B2(n[1967]), .ZN(
        n3949) );
  OAI221_X1 U1498 ( .B1(n570), .B2(n3222), .C1(n562), .C2(n3213), .A(n3953), 
        .ZN(n3952) );
  AOI22_X1 U1499 ( .A1(n3201), .A2(n[2087]), .B1(n3193), .B2(n[2095]), .ZN(
        n3953) );
  OAI221_X1 U1500 ( .B1(n2874), .B2(n3225), .C1(n2866), .C2(n3214), .A(n3861), 
        .ZN(n3860) );
  AOI22_X1 U1501 ( .A1(n3205), .A2(n[807]), .B1(n3191), .B2(n[815]), .ZN(n3861) );
  OAI221_X1 U1502 ( .B1(n2746), .B2(n3225), .C1(n2738), .C2(n3214), .A(n3865), 
        .ZN(n3864) );
  AOI22_X1 U1503 ( .A1(n3205), .A2(n[935]), .B1(n3194), .B2(n[943]), .ZN(n3865) );
  OAI221_X1 U1504 ( .B1(n2618), .B2(n3225), .C1(n2610), .C2(n3214), .A(n3869), 
        .ZN(n3868) );
  AOI22_X1 U1505 ( .A1(n3205), .A2(n[1063]), .B1(n3192), .B2(n[1071]), .ZN(
        n3869) );
  OAI221_X1 U1506 ( .B1(n2938), .B2(n3225), .C1(n2930), .C2(n3214), .A(n3881), 
        .ZN(n3880) );
  AOI22_X1 U1507 ( .A1(n3205), .A2(n[743]), .B1(n3190), .B2(n[751]), .ZN(n3881) );
  OAI221_X1 U1508 ( .B1(n2810), .B2(n3225), .C1(n2802), .C2(n3214), .A(n3885), 
        .ZN(n3884) );
  AOI22_X1 U1509 ( .A1(n3205), .A2(n[871]), .B1(n3196), .B2(n[879]), .ZN(n3885) );
  OAI221_X1 U1510 ( .B1(n2682), .B2(n3225), .C1(n2674), .C2(n3214), .A(n3889), 
        .ZN(n3888) );
  AOI22_X1 U1511 ( .A1(n3205), .A2(n[999]), .B1(n3671), .B2(n[1007]), .ZN(
        n3889) );
  OAI221_X1 U1512 ( .B1(n1721), .B2(n3224), .C1(n1713), .C2(n3216), .A(n3757), 
        .ZN(n3756) );
  AOI22_X1 U1513 ( .A1(n3207), .A2(n[1512]), .B1(n3190), .B2(n[1520]), .ZN(
        n3757) );
  OAI221_X1 U1514 ( .B1(n1081), .B2(n3226), .C1(n1073), .C2(n3215), .A(n3772), 
        .ZN(n3771) );
  AOI22_X1 U1515 ( .A1(n3206), .A2(n[1832]), .B1(n3197), .B2(n[1840]), .ZN(
        n3772) );
  OAI221_X1 U1516 ( .B1(n825), .B2(n3218), .C1(n817), .C2(n3215), .A(n3776), 
        .ZN(n3775) );
  AOI22_X1 U1517 ( .A1(n3206), .A2(n[1960]), .B1(n3671), .B2(n[1968]), .ZN(
        n3776) );
  OAI221_X1 U1518 ( .B1(n569), .B2(n3224), .C1(n561), .C2(n3215), .A(n3780), 
        .ZN(n3779) );
  AOI22_X1 U1519 ( .A1(n3206), .A2(n[2088]), .B1(n3671), .B2(n[2096]), .ZN(
        n3780) );
  OAI221_X1 U1520 ( .B1(n1209), .B2(n3221), .C1(n1201), .C2(n3215), .A(n3792), 
        .ZN(n3791) );
  AOI22_X1 U1521 ( .A1(n3206), .A2(n[1768]), .B1(n3671), .B2(n[1776]), .ZN(
        n3792) );
  OAI221_X1 U1522 ( .B1(n953), .B2(n3223), .C1(n945), .C2(n3215), .A(n3796), 
        .ZN(n3795) );
  AOI22_X1 U1523 ( .A1(n3206), .A2(n[1896]), .B1(n3671), .B2(n[1904]), .ZN(
        n3796) );
  OAI221_X1 U1524 ( .B1(n697), .B2(n3218), .C1(n689), .C2(n3215), .A(n3800), 
        .ZN(n3799) );
  AOI22_X1 U1525 ( .A1(n3206), .A2(n[2024]), .B1(n3671), .B2(n[2032]), .ZN(
        n3800) );
  OAI221_X1 U1526 ( .B1(n2937), .B2(n3219), .C1(n2929), .C2(n3216), .A(n3704), 
        .ZN(n3702) );
  AOI22_X1 U1527 ( .A1(n3207), .A2(n[744]), .B1(n3671), .B2(n[752]), .ZN(n3704) );
  OAI221_X1 U1528 ( .B1(n2809), .B2(n3224), .C1(n2801), .C2(n3216), .A(n3709), 
        .ZN(n3707) );
  AOI22_X1 U1529 ( .A1(n3207), .A2(n[872]), .B1(n3190), .B2(n[880]), .ZN(n3709) );
  OAI221_X1 U1530 ( .B1(n2681), .B2(n3222), .C1(n2673), .C2(n3216), .A(n3714), 
        .ZN(n3712) );
  AOI22_X1 U1531 ( .A1(n3207), .A2(n[1000]), .B1(n3190), .B2(n[1008]), .ZN(
        n3714) );
  OAI221_X1 U1532 ( .B1(n313), .B2(n3224), .C1(n305), .C2(n3215), .A(n3815), 
        .ZN(n3814) );
  AOI22_X1 U1533 ( .A1(n3206), .A2(n[2344]), .B1(n3671), .B2(n[2352]), .ZN(
        n3815) );
  OAI221_X1 U1534 ( .B1(n185), .B2(n3220), .C1(n177), .C2(n3215), .A(n3819), 
        .ZN(n3818) );
  AOI22_X1 U1535 ( .A1(n3206), .A2(n[2472]), .B1(n3671), .B2(n[2480]), .ZN(
        n3819) );
  OAI221_X1 U1536 ( .B1(n57), .B2(n3221), .C1(n49), .C2(n3215), .A(n3823), 
        .ZN(n3822) );
  AOI22_X1 U1537 ( .A1(n3206), .A2(n[2600]), .B1(n3671), .B2(n[2608]), .ZN(
        n3823) );
  OAI221_X1 U1538 ( .B1(n377), .B2(n3225), .C1(n369), .C2(n3214), .A(n3835), 
        .ZN(n3834) );
  AOI22_X1 U1539 ( .A1(n3205), .A2(n[2280]), .B1(n3195), .B2(n[2288]), .ZN(
        n3835) );
  OAI221_X1 U1540 ( .B1(n249), .B2(n3225), .C1(n241), .C2(n3214), .A(n3839), 
        .ZN(n3838) );
  AOI22_X1 U1541 ( .A1(n3205), .A2(n[2408]), .B1(n3193), .B2(n[2416]), .ZN(
        n3839) );
  OAI221_X1 U1542 ( .B1(n121), .B2(n3225), .C1(n113), .C2(n3214), .A(n3843), 
        .ZN(n3842) );
  AOI22_X1 U1543 ( .A1(n3205), .A2(n[2536]), .B1(n3196), .B2(n[2544]), .ZN(
        n3843) );
  AOI22_X1 U1544 ( .A1(n3670), .A2(n[675]), .B1(n3196), .B2(n[683]), .ZN(n4545) );
  AOI22_X1 U1545 ( .A1(n3205), .A2(n[803]), .B1(n3194), .B2(n[811]), .ZN(n4549) );
  AOI22_X1 U1546 ( .A1(n3202), .A2(n[931]), .B1(n3191), .B2(n[939]), .ZN(n4553) );
  AOI22_X1 U1547 ( .A1(n3207), .A2(n[1059]), .B1(n3192), .B2(n[1067]), .ZN(
        n4557) );
  AOI22_X1 U1548 ( .A1(n3206), .A2(n[611]), .B1(n3197), .B2(n[619]), .ZN(n4565) );
  AOI22_X1 U1549 ( .A1(n3200), .A2(n[739]), .B1(n3198), .B2(n[747]), .ZN(n4569) );
  AOI22_X1 U1550 ( .A1(n3199), .A2(n[867]), .B1(n3194), .B2(n[875]), .ZN(n4573) );
  AOI22_X1 U1551 ( .A1(n3670), .A2(n[1187]), .B1(n3191), .B2(n[1195]), .ZN(
        n4587) );
  AOI22_X1 U1552 ( .A1(n3207), .A2(n[1191]), .B1(n3190), .B2(n[1199]), .ZN(
        n3899) );
  AOI22_X1 U1553 ( .A1(n3670), .A2(n[1319]), .B1(n3192), .B2(n[1327]), .ZN(
        n3903) );
  AOI22_X1 U1554 ( .A1(n3203), .A2(n[1447]), .B1(n3192), .B2(n[1455]), .ZN(
        n3907) );
  AOI22_X1 U1555 ( .A1(n3205), .A2(n[1575]), .B1(n3192), .B2(n[1583]), .ZN(
        n3911) );
  AOI22_X1 U1556 ( .A1(n3202), .A2(n[1127]), .B1(n3195), .B2(n[1135]), .ZN(
        n3919) );
  AOI22_X1 U1557 ( .A1(n3207), .A2(n[1255]), .B1(n3192), .B2(n[1263]), .ZN(
        n3923) );
  AOI22_X1 U1558 ( .A1(n3204), .A2(n[1383]), .B1(n3191), .B2(n[1391]), .ZN(
        n3927) );
  AOI22_X1 U1559 ( .A1(n3201), .A2(n[1703]), .B1(n3198), .B2(n[1711]), .ZN(
        n3941) );
  OAI221_X1 U1560 ( .B1(n2841), .B2(n3182), .C1(n2833), .C2(n3180), .A(n3681), 
        .ZN(n3677) );
  AOI22_X1 U1561 ( .A1(n3171), .A2(n[776]), .B1(n3161), .B2(n[784]), .ZN(n3681) );
  OAI221_X1 U1562 ( .B1(n2713), .B2(n3187), .C1(n2705), .C2(n3180), .A(n3686), 
        .ZN(n3682) );
  AOI22_X1 U1563 ( .A1(n3171), .A2(n[904]), .B1(n3161), .B2(n[912]), .ZN(n3686) );
  OAI221_X1 U1564 ( .B1(n2553), .B2(n3188), .C1(n2545), .C2(n3180), .A(n3691), 
        .ZN(n3687) );
  AOI22_X1 U1565 ( .A1(n3171), .A2(n[1032]), .B1(n3161), .B2(n[1040]), .ZN(
        n3691) );
  OAI221_X1 U1566 ( .B1(n2654), .B2(n3185), .C1(n2646), .C2(n3673), .A(n4578), 
        .ZN(n4575) );
  AOI22_X1 U1567 ( .A1(n3675), .A2(n[963]), .B1(n3156), .B2(n[971]), .ZN(n4578) );
  OAI221_X1 U1568 ( .B1(n2046), .B2(n3184), .C1(n2038), .C2(n3180), .A(n4592), 
        .ZN(n4589) );
  AOI22_X1 U1569 ( .A1(n3164), .A2(n[1283]), .B1(n3157), .B2(n[1291]), .ZN(
        n4592) );
  OAI221_X1 U1570 ( .B1(n1790), .B2(n3184), .C1(n1782), .C2(n3180), .A(n4596), 
        .ZN(n4593) );
  AOI22_X1 U1571 ( .A1(n3169), .A2(n[1411]), .B1(n3154), .B2(n[1419]), .ZN(
        n4596) );
  OAI221_X1 U1572 ( .B1(n1534), .B2(n3189), .C1(n1526), .C2(n3180), .A(n4600), 
        .ZN(n4597) );
  AOI22_X1 U1573 ( .A1(n3168), .A2(n[1539]), .B1(n3160), .B2(n[1547]), .ZN(
        n4600) );
  OAI221_X1 U1574 ( .B1(n2653), .B2(n3672), .C1(n2645), .C2(n3177), .A(n4406), 
        .ZN(n4403) );
  AOI22_X1 U1575 ( .A1(n3168), .A2(n[964]), .B1(n3153), .B2(n[972]), .ZN(n4406) );
  OAI221_X1 U1576 ( .B1(n2045), .B2(n3181), .C1(n2037), .C2(n3175), .A(n4420), 
        .ZN(n4417) );
  AOI22_X1 U1577 ( .A1(n3675), .A2(n[1284]), .B1(n3161), .B2(n[1292]), .ZN(
        n4420) );
  OAI221_X1 U1578 ( .B1(n1789), .B2(n3185), .C1(n1781), .C2(n3177), .A(n4424), 
        .ZN(n4421) );
  AOI22_X1 U1579 ( .A1(n3162), .A2(n[1412]), .B1(n3161), .B2(n[1420]), .ZN(
        n4424) );
  OAI221_X1 U1580 ( .B1(n1533), .B2(n3186), .C1(n1525), .C2(n3178), .A(n4428), 
        .ZN(n4425) );
  AOI22_X1 U1581 ( .A1(n3171), .A2(n[1540]), .B1(n3156), .B2(n[1548]), .ZN(
        n4428) );
  OAI221_X1 U1582 ( .B1(n2173), .B2(n3183), .C1(n2165), .C2(n3174), .A(n4440), 
        .ZN(n4437) );
  AOI22_X1 U1583 ( .A1(n3163), .A2(n[1220]), .B1(n3161), .B2(n[1228]), .ZN(
        n4440) );
  OAI221_X1 U1584 ( .B1(n1917), .B2(n3187), .C1(n1909), .C2(n3177), .A(n4444), 
        .ZN(n4441) );
  AOI22_X1 U1585 ( .A1(n3168), .A2(n[1348]), .B1(n3156), .B2(n[1356]), .ZN(
        n4444) );
  OAI221_X1 U1586 ( .B1(n1661), .B2(n3185), .C1(n1653), .C2(n3176), .A(n4448), 
        .ZN(n4445) );
  AOI22_X1 U1587 ( .A1(n3165), .A2(n[1476]), .B1(n3676), .B2(n[1484]), .ZN(
        n4448) );
  OAI221_X1 U1588 ( .B1(n1021), .B2(n3185), .C1(n1013), .C2(n3174), .A(n4462), 
        .ZN(n4459) );
  AOI22_X1 U1589 ( .A1(n3169), .A2(n[1796]), .B1(n3161), .B2(n[1804]), .ZN(
        n4462) );
  OAI221_X1 U1590 ( .B1(n765), .B2(n3185), .C1(n757), .C2(n3179), .A(n4466), 
        .ZN(n4463) );
  AOI22_X1 U1591 ( .A1(n3170), .A2(n[1924]), .B1(n3159), .B2(n[1932]), .ZN(
        n4466) );
  OAI221_X1 U1592 ( .B1(n541), .B2(n3188), .C1(n533), .C2(n3180), .A(n4470), 
        .ZN(n4467) );
  AOI22_X1 U1593 ( .A1(n3167), .A2(n[2052]), .B1(n3161), .B2(n[2060]), .ZN(
        n4470) );
  OAI221_X1 U1594 ( .B1(n1149), .B2(n3188), .C1(n1141), .C2(n3178), .A(n4482), 
        .ZN(n4479) );
  AOI22_X1 U1595 ( .A1(n3171), .A2(n[1732]), .B1(n3161), .B2(n[1740]), .ZN(
        n4482) );
  OAI221_X1 U1596 ( .B1(n893), .B2(n3672), .C1(n885), .C2(n3175), .A(n4486), 
        .ZN(n4483) );
  AOI22_X1 U1597 ( .A1(n3171), .A2(n[1860]), .B1(n3160), .B2(n[1868]), .ZN(
        n4486) );
  OAI221_X1 U1598 ( .B1(n637), .B2(n3185), .C1(n629), .C2(n3173), .A(n4490), 
        .ZN(n4487) );
  AOI22_X1 U1599 ( .A1(n3167), .A2(n[1988]), .B1(n3161), .B2(n[1996]), .ZN(
        n4490) );
  OAI221_X1 U1600 ( .B1(n285), .B2(n3187), .C1(n277), .C2(n3174), .A(n4504), 
        .ZN(n4501) );
  AOI22_X1 U1601 ( .A1(n3171), .A2(n[2308]), .B1(n3158), .B2(n[2316]), .ZN(
        n4504) );
  OAI221_X1 U1602 ( .B1(n157), .B2(n3185), .C1(n149), .C2(n3178), .A(n4508), 
        .ZN(n4505) );
  AOI22_X1 U1603 ( .A1(n3171), .A2(n[2436]), .B1(n3158), .B2(n[2444]), .ZN(
        n4508) );
  OAI221_X1 U1604 ( .B1(n29), .B2(n3187), .C1(n21), .C2(n3172), .A(n4512), 
        .ZN(n4509) );
  AOI22_X1 U1605 ( .A1(n3171), .A2(n[2564]), .B1(n3159), .B2(n[2572]), .ZN(
        n4512) );
  OAI221_X1 U1606 ( .B1(n349), .B2(n3186), .C1(n341), .C2(n3175), .A(n4524), 
        .ZN(n4521) );
  AOI22_X1 U1607 ( .A1(n3171), .A2(n[2244]), .B1(n3155), .B2(n[2252]), .ZN(
        n4524) );
  OAI221_X1 U1608 ( .B1(n221), .B2(n3184), .C1(n213), .C2(n3177), .A(n4528), 
        .ZN(n4525) );
  AOI22_X1 U1609 ( .A1(n3167), .A2(n[2372]), .B1(n3157), .B2(n[2380]), .ZN(
        n4528) );
  OAI221_X1 U1610 ( .B1(n93), .B2(n3187), .C1(n85), .C2(n3178), .A(n4532), 
        .ZN(n4529) );
  AOI22_X1 U1611 ( .A1(n3164), .A2(n[2500]), .B1(n3156), .B2(n[2508]), .ZN(
        n4532) );
  OAI221_X1 U1612 ( .B1(n348), .B2(n3183), .C1(n340), .C2(n3673), .A(n4352), 
        .ZN(n4349) );
  AOI22_X1 U1613 ( .A1(n3163), .A2(n[2245]), .B1(n3676), .B2(n[2253]), .ZN(
        n4352) );
  OAI221_X1 U1614 ( .B1(n220), .B2(n3183), .C1(n212), .C2(n3172), .A(n4356), 
        .ZN(n4353) );
  AOI22_X1 U1615 ( .A1(n3169), .A2(n[2373]), .B1(n3158), .B2(n[2381]), .ZN(
        n4356) );
  OAI221_X1 U1616 ( .B1(n92), .B2(n3182), .C1(n84), .C2(n3179), .A(n4360), 
        .ZN(n4357) );
  AOI22_X1 U1617 ( .A1(n3171), .A2(n[2501]), .B1(n3154), .B2(n[2509]), .ZN(
        n4360) );
  OAI221_X1 U1618 ( .B1(n1658), .B2(n3181), .C1(n1650), .C2(n3176), .A(n3932), 
        .ZN(n3929) );
  AOI22_X1 U1619 ( .A1(n3675), .A2(n[1479]), .B1(n3157), .B2(n[1487]), .ZN(
        n3932) );
  OAI221_X1 U1620 ( .B1(n1018), .B2(n3181), .C1(n1010), .C2(n3176), .A(n3946), 
        .ZN(n3943) );
  AOI22_X1 U1621 ( .A1(n3164), .A2(n[1799]), .B1(n3157), .B2(n[1807]), .ZN(
        n3946) );
  OAI221_X1 U1622 ( .B1(n762), .B2(n3181), .C1(n754), .C2(n3176), .A(n3950), 
        .ZN(n3947) );
  AOI22_X1 U1623 ( .A1(n3166), .A2(n[1927]), .B1(n3157), .B2(n[1935]), .ZN(
        n3950) );
  OAI221_X1 U1624 ( .B1(n538), .B2(n3181), .C1(n530), .C2(n3176), .A(n3954), 
        .ZN(n3951) );
  AOI22_X1 U1625 ( .A1(n3170), .A2(n[2055]), .B1(n3157), .B2(n[2063]), .ZN(
        n3954) );
  OAI221_X1 U1626 ( .B1(n2842), .B2(n3181), .C1(n2834), .C2(n3177), .A(n3862), 
        .ZN(n3859) );
  AOI22_X1 U1627 ( .A1(n3168), .A2(n[775]), .B1(n3158), .B2(n[783]), .ZN(n3862) );
  OAI221_X1 U1628 ( .B1(n2714), .B2(n3187), .C1(n2706), .C2(n3177), .A(n3866), 
        .ZN(n3863) );
  AOI22_X1 U1629 ( .A1(n3168), .A2(n[903]), .B1(n3158), .B2(n[911]), .ZN(n3866) );
  OAI221_X1 U1630 ( .B1(n2554), .B2(n3182), .C1(n2546), .C2(n3177), .A(n3870), 
        .ZN(n3867) );
  AOI22_X1 U1631 ( .A1(n3168), .A2(n[1031]), .B1(n3158), .B2(n[1039]), .ZN(
        n3870) );
  OAI221_X1 U1632 ( .B1(n2906), .B2(n3182), .C1(n2898), .C2(n3177), .A(n3882), 
        .ZN(n3879) );
  AOI22_X1 U1633 ( .A1(n3168), .A2(n[711]), .B1(n3158), .B2(n[719]), .ZN(n3882) );
  OAI221_X1 U1634 ( .B1(n2778), .B2(n3183), .C1(n2770), .C2(n3177), .A(n3886), 
        .ZN(n3883) );
  AOI22_X1 U1635 ( .A1(n3168), .A2(n[839]), .B1(n3158), .B2(n[847]), .ZN(n3886) );
  OAI221_X1 U1636 ( .B1(n2650), .B2(n3184), .C1(n2642), .C2(n3177), .A(n3890), 
        .ZN(n3887) );
  AOI22_X1 U1637 ( .A1(n3168), .A2(n[967]), .B1(n3158), .B2(n[975]), .ZN(n3890) );
  OAI221_X1 U1638 ( .B1(n1657), .B2(n3672), .C1(n1649), .C2(n3179), .A(n3758), 
        .ZN(n3755) );
  AOI22_X1 U1639 ( .A1(n3170), .A2(n[1480]), .B1(n3160), .B2(n[1488]), .ZN(
        n3758) );
  OAI221_X1 U1640 ( .B1(n1017), .B2(n3188), .C1(n1009), .C2(n3178), .A(n3773), 
        .ZN(n3770) );
  AOI22_X1 U1641 ( .A1(n3169), .A2(n[1800]), .B1(n3159), .B2(n[1808]), .ZN(
        n3773) );
  OAI221_X1 U1642 ( .B1(n761), .B2(n3188), .C1(n753), .C2(n3178), .A(n3777), 
        .ZN(n3774) );
  AOI22_X1 U1643 ( .A1(n3169), .A2(n[1928]), .B1(n3159), .B2(n[1936]), .ZN(
        n3777) );
  OAI221_X1 U1644 ( .B1(n537), .B2(n3189), .C1(n529), .C2(n3178), .A(n3781), 
        .ZN(n3778) );
  AOI22_X1 U1645 ( .A1(n3169), .A2(n[2056]), .B1(n3159), .B2(n[2064]), .ZN(
        n3781) );
  OAI221_X1 U1646 ( .B1(n1145), .B2(n3182), .C1(n1137), .C2(n3178), .A(n3793), 
        .ZN(n3790) );
  AOI22_X1 U1647 ( .A1(n3169), .A2(n[1736]), .B1(n3159), .B2(n[1744]), .ZN(
        n3793) );
  OAI221_X1 U1648 ( .B1(n889), .B2(n3183), .C1(n881), .C2(n3178), .A(n3797), 
        .ZN(n3794) );
  AOI22_X1 U1649 ( .A1(n3169), .A2(n[1864]), .B1(n3159), .B2(n[1872]), .ZN(
        n3797) );
  OAI221_X1 U1650 ( .B1(n633), .B2(n3189), .C1(n625), .C2(n3178), .A(n3801), 
        .ZN(n3798) );
  AOI22_X1 U1651 ( .A1(n3169), .A2(n[1992]), .B1(n3159), .B2(n[2000]), .ZN(
        n3801) );
  OAI221_X1 U1652 ( .B1(n2905), .B2(n3186), .C1(n2897), .C2(n3179), .A(n3705), 
        .ZN(n3701) );
  AOI22_X1 U1653 ( .A1(n3170), .A2(n[712]), .B1(n3160), .B2(n[720]), .ZN(n3705) );
  OAI221_X1 U1654 ( .B1(n2777), .B2(n3672), .C1(n2769), .C2(n3179), .A(n3710), 
        .ZN(n3706) );
  AOI22_X1 U1655 ( .A1(n3170), .A2(n[840]), .B1(n3160), .B2(n[848]), .ZN(n3710) );
  OAI221_X1 U1656 ( .B1(n2649), .B2(n3672), .C1(n2641), .C2(n3179), .A(n3715), 
        .ZN(n3711) );
  AOI22_X1 U1657 ( .A1(n3170), .A2(n[968]), .B1(n3160), .B2(n[976]), .ZN(n3715) );
  OAI221_X1 U1658 ( .B1(n281), .B2(n3186), .C1(n273), .C2(n3178), .A(n3816), 
        .ZN(n3813) );
  AOI22_X1 U1659 ( .A1(n3169), .A2(n[2312]), .B1(n3159), .B2(n[2320]), .ZN(
        n3816) );
  OAI221_X1 U1660 ( .B1(n153), .B2(n3182), .C1(n145), .C2(n3178), .A(n3820), 
        .ZN(n3817) );
  AOI22_X1 U1661 ( .A1(n3169), .A2(n[2440]), .B1(n3159), .B2(n[2448]), .ZN(
        n3820) );
  OAI221_X1 U1662 ( .B1(n25), .B2(n3181), .C1(n17), .C2(n3178), .A(n3824), 
        .ZN(n3821) );
  AOI22_X1 U1663 ( .A1(n3169), .A2(n[2568]), .B1(n3159), .B2(n[2576]), .ZN(
        n3824) );
  OAI221_X1 U1664 ( .B1(n345), .B2(n3182), .C1(n337), .C2(n3177), .A(n3836), 
        .ZN(n3833) );
  AOI22_X1 U1665 ( .A1(n3168), .A2(n[2248]), .B1(n3158), .B2(n[2256]), .ZN(
        n3836) );
  OAI221_X1 U1666 ( .B1(n217), .B2(n3183), .C1(n209), .C2(n3177), .A(n3840), 
        .ZN(n3837) );
  AOI22_X1 U1667 ( .A1(n3168), .A2(n[2376]), .B1(n3158), .B2(n[2384]), .ZN(
        n3840) );
  OAI221_X1 U1668 ( .B1(n89), .B2(n3188), .C1(n81), .C2(n3177), .A(n3844), 
        .ZN(n3841) );
  AOI22_X1 U1669 ( .A1(n3168), .A2(n[2504]), .B1(n3158), .B2(n[2512]), .ZN(
        n3844) );
  AOI22_X1 U1670 ( .A1(n3205), .A2(n[676]), .B1(n3671), .B2(n[684]), .ZN(n4373) );
  AOI22_X1 U1671 ( .A1(n3199), .A2(n[804]), .B1(n3193), .B2(n[812]), .ZN(n4377) );
  AOI22_X1 U1672 ( .A1(n3204), .A2(n[932]), .B1(n3195), .B2(n[940]), .ZN(n4381) );
  AOI22_X1 U1673 ( .A1(n3204), .A2(n[1060]), .B1(n3195), .B2(n[1068]), .ZN(
        n4385) );
  AOI22_X1 U1674 ( .A1(n3206), .A2(n[612]), .B1(n3671), .B2(n[620]), .ZN(n4393) );
  AOI22_X1 U1675 ( .A1(n3203), .A2(n[740]), .B1(n3197), .B2(n[748]), .ZN(n4397) );
  AOI22_X1 U1676 ( .A1(n3199), .A2(n[868]), .B1(n3193), .B2(n[876]), .ZN(n4401) );
  AOI22_X1 U1677 ( .A1(n3670), .A2(n[1188]), .B1(n3198), .B2(n[1196]), .ZN(
        n4415) );
  AOI22_X1 U1678 ( .A1(n3207), .A2(n[1124]), .B1(n3191), .B2(n[1132]), .ZN(
        n4435) );
  AOI22_X1 U1679 ( .A1(n3206), .A2(n[1700]), .B1(n3196), .B2(n[1708]), .ZN(
        n4457) );
  AOI22_X1 U1680 ( .A1(n3208), .A2(n[1636]), .B1(n3191), .B2(n[1644]), .ZN(
        n4477) );
  AOI22_X1 U1681 ( .A1(n3208), .A2(n[2212]), .B1(n3198), .B2(n[2220]), .ZN(
        n4499) );
  AOI22_X1 U1682 ( .A1(n3208), .A2(n[2148]), .B1(n3192), .B2(n[2156]), .ZN(
        n4519) );
  AOI22_X1 U1683 ( .A1(n3206), .A2(n[2149]), .B1(n3196), .B2(n[2157]), .ZN(
        n4347) );
  AOI22_X1 U1684 ( .A1(n3205), .A2(n[679]), .B1(n3192), .B2(n[687]), .ZN(n3857) );
  AOI22_X1 U1685 ( .A1(n3205), .A2(n[615]), .B1(n3192), .B2(n[623]), .ZN(n3877) );
  AOI22_X1 U1686 ( .A1(n3207), .A2(n[1192]), .B1(n3195), .B2(n[1200]), .ZN(
        n3725) );
  AOI22_X1 U1687 ( .A1(n3207), .A2(n[1320]), .B1(n3196), .B2(n[1328]), .ZN(
        n3729) );
  AOI22_X1 U1688 ( .A1(n3207), .A2(n[1448]), .B1(n3671), .B2(n[1456]), .ZN(
        n3733) );
  AOI22_X1 U1689 ( .A1(n3207), .A2(n[1576]), .B1(n3190), .B2(n[1584]), .ZN(
        n3737) );
  AOI22_X1 U1690 ( .A1(n3207), .A2(n[1128]), .B1(n3671), .B2(n[1136]), .ZN(
        n3745) );
  AOI22_X1 U1691 ( .A1(n3207), .A2(n[1256]), .B1(n3193), .B2(n[1264]), .ZN(
        n3749) );
  AOI22_X1 U1692 ( .A1(n3207), .A2(n[1384]), .B1(n3190), .B2(n[1392]), .ZN(
        n3753) );
  AOI22_X1 U1693 ( .A1(n3206), .A2(n[1704]), .B1(n3671), .B2(n[1712]), .ZN(
        n3768) );
  AOI22_X1 U1694 ( .A1(n3206), .A2(n[1640]), .B1(n3671), .B2(n[1648]), .ZN(
        n3788) );
  AOI22_X1 U1695 ( .A1(n3207), .A2(n[616]), .B1(n3194), .B2(n[624]), .ZN(n3699) );
  AOI22_X1 U1696 ( .A1(n3208), .A2(n[680]), .B1(n3190), .B2(n[688]), .ZN(n3669) );
  AOI22_X1 U1697 ( .A1(n3206), .A2(n[2216]), .B1(n3671), .B2(n[2224]), .ZN(
        n3811) );
  AOI22_X1 U1698 ( .A1(n3205), .A2(n[2152]), .B1(n3198), .B2(n[2160]), .ZN(
        n3831) );
  OAI22_X1 U1699 ( .A1(n3350), .A2(n3145), .B1(n3296), .B2(n1952), .ZN(n5840)
         );
  OAI22_X1 U1700 ( .A1(n3350), .A2(n3128), .B1(n3296), .B2(n1951), .ZN(n5841)
         );
  OAI22_X1 U1701 ( .A1(n3350), .A2(n7256), .B1(n3296), .B2(n1950), .ZN(n5842)
         );
  OAI22_X1 U1702 ( .A1(n3349), .A2(n3145), .B1(n7117), .B2(n1976), .ZN(n5832)
         );
  OAI22_X1 U1703 ( .A1(n3349), .A2(n3130), .B1(n7117), .B2(n1975), .ZN(n5833)
         );
  OAI22_X1 U1704 ( .A1(n3349), .A2(n7256), .B1(n7117), .B2(n1974), .ZN(n5834)
         );
  OAI22_X1 U1705 ( .A1(n3349), .A2(n7255), .B1(n7117), .B2(n1973), .ZN(n5835)
         );
  OAI22_X1 U1706 ( .A1(n3349), .A2(n3106), .B1(n7117), .B2(n1972), .ZN(n5836)
         );
  OAI22_X1 U1707 ( .A1(n3349), .A2(n3091), .B1(n7117), .B2(n1971), .ZN(n5837)
         );
  OAI22_X1 U1708 ( .A1(n3349), .A2(n3083), .B1(n7117), .B2(n1970), .ZN(n5838)
         );
  OAI22_X1 U1709 ( .A1(n3349), .A2(n3074), .B1(n7117), .B2(n1969), .ZN(n5839)
         );
  OAI21_X1 U1710 ( .B1(n4887), .B2(n4888), .A(n3227), .ZN(n4886) );
  OAI221_X1 U1711 ( .B1(n2976), .B2(n3672), .C1(n2968), .C2(n3180), .A(n4890), 
        .ZN(n4887) );
  OAI221_X1 U1712 ( .B1(n3008), .B2(n3225), .C1(n3000), .C2(n3209), .A(n4889), 
        .ZN(n4888) );
  AOI22_X1 U1713 ( .A1(n3675), .A2(n[641]), .B1(n3153), .B2(n[649]), .ZN(n4890) );
  OAI21_X1 U1714 ( .B1(n4907), .B2(n4908), .A(n3149), .ZN(n4906) );
  OAI221_X1 U1715 ( .B1(n3040), .B2(n3185), .C1(n3032), .C2(n3673), .A(n4910), 
        .ZN(n4907) );
  OAI221_X1 U1716 ( .B1(n3072), .B2(n3218), .C1(n3064), .C2(n3668), .A(n4909), 
        .ZN(n4908) );
  AOI22_X1 U1717 ( .A1(n3163), .A2(n[577]), .B1(n3160), .B2(n[585]), .ZN(n4910) );
  OAI21_X1 U1718 ( .B1(n4929), .B2(n4930), .A(n3227), .ZN(n4928) );
  OAI221_X1 U1719 ( .B1(n2304), .B2(n3184), .C1(n2296), .C2(n3178), .A(n4932), 
        .ZN(n4929) );
  OAI221_X1 U1720 ( .B1(n2368), .B2(n3226), .C1(n2360), .C2(n3209), .A(n4931), 
        .ZN(n4930) );
  AOI22_X1 U1721 ( .A1(n3171), .A2(n[1153]), .B1(n3676), .B2(n[1161]), .ZN(
        n4932) );
  OAI21_X1 U1722 ( .B1(n4949), .B2(n4950), .A(n3149), .ZN(n4948) );
  OAI221_X1 U1723 ( .B1(n2432), .B2(n3186), .C1(n2424), .C2(n3172), .A(n4952), 
        .ZN(n4949) );
  OAI221_X1 U1724 ( .B1(n2496), .B2(n3225), .C1(n2488), .C2(n3209), .A(n4951), 
        .ZN(n4950) );
  AOI22_X1 U1725 ( .A1(n3168), .A2(n[1089]), .B1(n3156), .B2(n[1097]), .ZN(
        n4952) );
  OAI21_X1 U1726 ( .B1(n4971), .B2(n4972), .A(n3227), .ZN(n4970) );
  OAI221_X1 U1727 ( .B1(n1280), .B2(n3189), .C1(n1272), .C2(n3172), .A(n4974), 
        .ZN(n4971) );
  OAI221_X1 U1728 ( .B1(n1344), .B2(n3222), .C1(n1336), .C2(n3210), .A(n4973), 
        .ZN(n4972) );
  AOI22_X1 U1729 ( .A1(n3166), .A2(n[1665]), .B1(n3161), .B2(n[1673]), .ZN(
        n4974) );
  OAI21_X1 U1730 ( .B1(n4991), .B2(n4992), .A(n3149), .ZN(n4990) );
  OAI221_X1 U1731 ( .B1(n1408), .B2(n3182), .C1(n1400), .C2(n3174), .A(n4994), 
        .ZN(n4991) );
  OAI221_X1 U1732 ( .B1(n1472), .B2(n3221), .C1(n1464), .C2(n3210), .A(n4993), 
        .ZN(n4992) );
  AOI22_X1 U1733 ( .A1(n3167), .A2(n[1601]), .B1(n3158), .B2(n[1609]), .ZN(
        n4994) );
  OAI21_X1 U1734 ( .B1(n5013), .B2(n5014), .A(n3227), .ZN(n5012) );
  OAI221_X1 U1735 ( .B1(n416), .B2(n3182), .C1(n408), .C2(n3175), .A(n5017), 
        .ZN(n5013) );
  OAI221_X1 U1736 ( .B1(n448), .B2(n3225), .C1(n440), .C2(n3215), .A(n5016), 
        .ZN(n5014) );
  AOI22_X1 U1737 ( .A1(n3163), .A2(n[2177]), .B1(n3154), .B2(n[2185]), .ZN(
        n5017) );
  OAI21_X1 U1738 ( .B1(n5037), .B2(n5038), .A(n3149), .ZN(n5036) );
  OAI221_X1 U1739 ( .B1(n480), .B2(n3182), .C1(n472), .C2(n3178), .A(n5040), 
        .ZN(n5037) );
  OAI221_X1 U1740 ( .B1(n512), .B2(n3667), .C1(n504), .C2(n3216), .A(n5039), 
        .ZN(n5038) );
  AOI22_X1 U1741 ( .A1(n3168), .A2(n[2113]), .B1(n3156), .B2(n[2121]), .ZN(
        n5040) );
  OAI21_X1 U1742 ( .B1(n4715), .B2(n4716), .A(n3227), .ZN(n4714) );
  OAI221_X1 U1743 ( .B1(n2975), .B2(n3181), .C1(n2967), .C2(n3172), .A(n4718), 
        .ZN(n4715) );
  OAI221_X1 U1744 ( .B1(n3007), .B2(n3218), .C1(n2999), .C2(n3213), .A(n4717), 
        .ZN(n4716) );
  AOI22_X1 U1745 ( .A1(n3168), .A2(n[642]), .B1(n3159), .B2(n[650]), .ZN(n4718) );
  OAI21_X1 U1746 ( .B1(n4735), .B2(n4736), .A(n3149), .ZN(n4734) );
  OAI221_X1 U1747 ( .B1(n3039), .B2(n3182), .C1(n3031), .C2(n3180), .A(n4738), 
        .ZN(n4735) );
  OAI221_X1 U1748 ( .B1(n3071), .B2(n3220), .C1(n3063), .C2(n3668), .A(n4737), 
        .ZN(n4736) );
  AOI22_X1 U1749 ( .A1(n3168), .A2(n[578]), .B1(n3153), .B2(n[586]), .ZN(n4738) );
  OAI21_X1 U1750 ( .B1(n4757), .B2(n4758), .A(n3227), .ZN(n4756) );
  OAI221_X1 U1751 ( .B1(n2303), .B2(n3183), .C1(n2295), .C2(n3673), .A(n4760), 
        .ZN(n4757) );
  OAI221_X1 U1752 ( .B1(n2367), .B2(n3225), .C1(n2359), .C2(n3668), .A(n4759), 
        .ZN(n4758) );
  AOI22_X1 U1753 ( .A1(n3169), .A2(n[1154]), .B1(n3159), .B2(n[1162]), .ZN(
        n4760) );
  OAI21_X1 U1754 ( .B1(n4777), .B2(n4778), .A(n3149), .ZN(n4776) );
  OAI221_X1 U1755 ( .B1(n2431), .B2(n3189), .C1(n2423), .C2(n3175), .A(n4780), 
        .ZN(n4777) );
  OAI221_X1 U1756 ( .B1(n2495), .B2(n3224), .C1(n2487), .C2(n3209), .A(n4779), 
        .ZN(n4778) );
  AOI22_X1 U1757 ( .A1(n3170), .A2(n[1090]), .B1(n3154), .B2(n[1098]), .ZN(
        n4780) );
  OAI21_X1 U1758 ( .B1(n4799), .B2(n4800), .A(n3227), .ZN(n4798) );
  OAI221_X1 U1759 ( .B1(n1279), .B2(n3183), .C1(n1271), .C2(n3174), .A(n4802), 
        .ZN(n4799) );
  OAI221_X1 U1760 ( .B1(n1343), .B2(n3223), .C1(n1335), .C2(n3211), .A(n4801), 
        .ZN(n4800) );
  AOI22_X1 U1761 ( .A1(n3170), .A2(n[1666]), .B1(n3676), .B2(n[1674]), .ZN(
        n4802) );
  OAI21_X1 U1762 ( .B1(n4819), .B2(n4820), .A(n3149), .ZN(n4818) );
  OAI221_X1 U1763 ( .B1(n1407), .B2(n3183), .C1(n1399), .C2(n3179), .A(n4822), 
        .ZN(n4819) );
  OAI221_X1 U1764 ( .B1(n1471), .B2(n3222), .C1(n1463), .C2(n3212), .A(n4821), 
        .ZN(n4820) );
  AOI22_X1 U1765 ( .A1(n3166), .A2(n[1602]), .B1(n3676), .B2(n[1610]), .ZN(
        n4822) );
  OAI21_X1 U1766 ( .B1(n4841), .B2(n4842), .A(n3227), .ZN(n4840) );
  OAI221_X1 U1767 ( .B1(n415), .B2(n3183), .C1(n407), .C2(n3172), .A(n4844), 
        .ZN(n4841) );
  OAI221_X1 U1768 ( .B1(n447), .B2(n3225), .C1(n439), .C2(n3209), .A(n4843), 
        .ZN(n4842) );
  AOI22_X1 U1769 ( .A1(n3170), .A2(n[2178]), .B1(n3676), .B2(n[2186]), .ZN(
        n4844) );
  OAI21_X1 U1770 ( .B1(n4861), .B2(n4862), .A(n3149), .ZN(n4860) );
  OAI221_X1 U1771 ( .B1(n479), .B2(n3188), .C1(n471), .C2(n3673), .A(n4864), 
        .ZN(n4861) );
  OAI221_X1 U1772 ( .B1(n511), .B2(n3223), .C1(n503), .C2(n3668), .A(n4863), 
        .ZN(n4862) );
  AOI22_X1 U1773 ( .A1(n3169), .A2(n[2114]), .B1(n3153), .B2(n[2122]), .ZN(
        n4864) );
  OAI21_X1 U1774 ( .B1(n4627), .B2(n4628), .A(n3666), .ZN(n4626) );
  OAI221_X1 U1775 ( .B1(n1278), .B2(n3183), .C1(n1270), .C2(n3173), .A(n4630), 
        .ZN(n4627) );
  OAI221_X1 U1776 ( .B1(n1342), .B2(n3226), .C1(n1334), .C2(n3668), .A(n4629), 
        .ZN(n4628) );
  AOI22_X1 U1777 ( .A1(n3166), .A2(n[1667]), .B1(n3157), .B2(n[1675]), .ZN(
        n4630) );
  OAI21_X1 U1778 ( .B1(n4647), .B2(n4648), .A(n3698), .ZN(n4646) );
  OAI221_X1 U1779 ( .B1(n1406), .B2(n3187), .C1(n1398), .C2(n3177), .A(n4650), 
        .ZN(n4647) );
  OAI221_X1 U1780 ( .B1(n1470), .B2(n3226), .C1(n1462), .C2(n3668), .A(n4649), 
        .ZN(n4648) );
  AOI22_X1 U1781 ( .A1(n3163), .A2(n[1603]), .B1(n3159), .B2(n[1611]), .ZN(
        n4650) );
  OAI21_X1 U1782 ( .B1(n4605), .B2(n4606), .A(n3698), .ZN(n4604) );
  OAI221_X1 U1783 ( .B1(n2430), .B2(n3184), .C1(n2422), .C2(n3178), .A(n4608), 
        .ZN(n4605) );
  OAI221_X1 U1784 ( .B1(n2494), .B2(n3226), .C1(n2486), .C2(n3209), .A(n4607), 
        .ZN(n4606) );
  AOI22_X1 U1785 ( .A1(n3675), .A2(n[1091]), .B1(n3160), .B2(n[1099]), .ZN(
        n4608) );
  OAI21_X1 U1786 ( .B1(n4669), .B2(n4670), .A(n3666), .ZN(n4668) );
  OAI221_X1 U1787 ( .B1(n414), .B2(n3182), .C1(n406), .C2(n3177), .A(n4672), 
        .ZN(n4669) );
  OAI221_X1 U1788 ( .B1(n446), .B2(n3218), .C1(n438), .C2(n3211), .A(n4671), 
        .ZN(n4670) );
  AOI22_X1 U1789 ( .A1(n3162), .A2(n[2179]), .B1(n3158), .B2(n[2187]), .ZN(
        n4672) );
  OAI21_X1 U1790 ( .B1(n4689), .B2(n4690), .A(n3698), .ZN(n4688) );
  OAI221_X1 U1791 ( .B1(n478), .B2(n3181), .C1(n470), .C2(n3673), .A(n4692), 
        .ZN(n4689) );
  OAI221_X1 U1792 ( .B1(n510), .B2(n3218), .C1(n502), .C2(n3668), .A(n4691), 
        .ZN(n4690) );
  AOI22_X1 U1793 ( .A1(n3170), .A2(n[2115]), .B1(n3159), .B2(n[2123]), .ZN(
        n4692) );
  OAI21_X1 U1794 ( .B1(n4199), .B2(n4200), .A(n3666), .ZN(n4198) );
  OAI221_X1 U1795 ( .B1(n2972), .B2(n3186), .C1(n2964), .C2(n3176), .A(n4202), 
        .ZN(n4199) );
  OAI221_X1 U1796 ( .B1(n3004), .B2(n3221), .C1(n2996), .C2(n3217), .A(n4201), 
        .ZN(n4200) );
  AOI22_X1 U1797 ( .A1(n3164), .A2(n[645]), .B1(n3159), .B2(n[653]), .ZN(n4202) );
  OAI21_X1 U1798 ( .B1(n4219), .B2(n4220), .A(n3698), .ZN(n4218) );
  OAI221_X1 U1799 ( .B1(n3036), .B2(n3185), .C1(n3028), .C2(n3174), .A(n4222), 
        .ZN(n4219) );
  OAI221_X1 U1800 ( .B1(n3068), .B2(n3220), .C1(n3060), .C2(n3211), .A(n4221), 
        .ZN(n4220) );
  AOI22_X1 U1801 ( .A1(n3163), .A2(n[581]), .B1(n3155), .B2(n[589]), .ZN(n4222) );
  OAI21_X1 U1802 ( .B1(n4241), .B2(n4242), .A(n3666), .ZN(n4240) );
  OAI221_X1 U1803 ( .B1(n2300), .B2(n3185), .C1(n2292), .C2(n3174), .A(n4244), 
        .ZN(n4241) );
  OAI221_X1 U1804 ( .B1(n2364), .B2(n3220), .C1(n2356), .C2(n3211), .A(n4243), 
        .ZN(n4242) );
  AOI22_X1 U1805 ( .A1(n3163), .A2(n[1157]), .B1(n3155), .B2(n[1165]), .ZN(
        n4244) );
  OAI21_X1 U1806 ( .B1(n4261), .B2(n4262), .A(n3698), .ZN(n4260) );
  OAI221_X1 U1807 ( .B1(n2428), .B2(n3185), .C1(n2420), .C2(n3174), .A(n4264), 
        .ZN(n4261) );
  OAI221_X1 U1808 ( .B1(n2492), .B2(n3220), .C1(n2484), .C2(n3211), .A(n4263), 
        .ZN(n4262) );
  AOI22_X1 U1809 ( .A1(n3163), .A2(n[1093]), .B1(n3155), .B2(n[1101]), .ZN(
        n4264) );
  OAI21_X1 U1810 ( .B1(n4283), .B2(n4284), .A(n3666), .ZN(n4282) );
  OAI221_X1 U1811 ( .B1(n1276), .B2(n3184), .C1(n1268), .C2(n3173), .A(n4286), 
        .ZN(n4283) );
  OAI221_X1 U1812 ( .B1(n1340), .B2(n3219), .C1(n1332), .C2(n3210), .A(n4285), 
        .ZN(n4284) );
  AOI22_X1 U1813 ( .A1(n3162), .A2(n[1669]), .B1(n3154), .B2(n[1677]), .ZN(
        n4286) );
  OAI21_X1 U1814 ( .B1(n4303), .B2(n4304), .A(n3698), .ZN(n4302) );
  OAI221_X1 U1815 ( .B1(n1404), .B2(n3184), .C1(n1396), .C2(n3173), .A(n4306), 
        .ZN(n4303) );
  OAI221_X1 U1816 ( .B1(n1468), .B2(n3219), .C1(n1460), .C2(n3210), .A(n4305), 
        .ZN(n4304) );
  AOI22_X1 U1817 ( .A1(n3162), .A2(n[1605]), .B1(n3154), .B2(n[1613]), .ZN(
        n4306) );
  OAI21_X1 U1818 ( .B1(n4325), .B2(n4326), .A(n3666), .ZN(n4324) );
  OAI221_X1 U1819 ( .B1(n412), .B2(n3184), .C1(n404), .C2(n3173), .A(n4328), 
        .ZN(n4325) );
  OAI221_X1 U1820 ( .B1(n444), .B2(n3219), .C1(n436), .C2(n3210), .A(n4327), 
        .ZN(n4326) );
  AOI22_X1 U1821 ( .A1(n3162), .A2(n[2181]), .B1(n3154), .B2(n[2189]), .ZN(
        n4328) );
  OAI21_X1 U1822 ( .B1(n4027), .B2(n4028), .A(n3227), .ZN(n4026) );
  OAI221_X1 U1823 ( .B1(n2971), .B2(n3188), .C1(n2963), .C2(n3178), .A(n4030), 
        .ZN(n4027) );
  OAI221_X1 U1824 ( .B1(n3003), .B2(n3223), .C1(n2995), .C2(n3213), .A(n4029), 
        .ZN(n4028) );
  AOI22_X1 U1825 ( .A1(n3166), .A2(n[646]), .B1(n3155), .B2(n[654]), .ZN(n4030) );
  OAI21_X1 U1826 ( .B1(n4047), .B2(n4048), .A(n3149), .ZN(n4046) );
  OAI221_X1 U1827 ( .B1(n3035), .B2(n3188), .C1(n3027), .C2(n3172), .A(n4050), 
        .ZN(n4047) );
  OAI221_X1 U1828 ( .B1(n3067), .B2(n3223), .C1(n3059), .C2(n3216), .A(n4049), 
        .ZN(n4048) );
  AOI22_X1 U1829 ( .A1(n3166), .A2(n[582]), .B1(n3155), .B2(n[590]), .ZN(n4050) );
  OAI21_X1 U1830 ( .B1(n4069), .B2(n4070), .A(n3227), .ZN(n4068) );
  OAI221_X1 U1831 ( .B1(n2299), .B2(n3188), .C1(n2291), .C2(n3179), .A(n4072), 
        .ZN(n4069) );
  OAI221_X1 U1832 ( .B1(n2363), .B2(n3223), .C1(n2355), .C2(n3215), .A(n4071), 
        .ZN(n4070) );
  AOI22_X1 U1833 ( .A1(n3166), .A2(n[1158]), .B1(n3160), .B2(n[1166]), .ZN(
        n4072) );
  OAI21_X1 U1834 ( .B1(n4089), .B2(n4090), .A(n3149), .ZN(n4088) );
  OAI221_X1 U1835 ( .B1(n2427), .B2(n3187), .C1(n2419), .C2(n3179), .A(n4092), 
        .ZN(n4089) );
  OAI221_X1 U1836 ( .B1(n2491), .B2(n3222), .C1(n2483), .C2(n3213), .A(n4091), 
        .ZN(n4090) );
  AOI22_X1 U1837 ( .A1(n3165), .A2(n[1094]), .B1(n3156), .B2(n[1102]), .ZN(
        n4092) );
  OAI21_X1 U1838 ( .B1(n4111), .B2(n4112), .A(n3666), .ZN(n4110) );
  OAI221_X1 U1839 ( .B1(n1275), .B2(n3187), .C1(n1267), .C2(n3174), .A(n4114), 
        .ZN(n4111) );
  OAI221_X1 U1840 ( .B1(n1339), .B2(n3222), .C1(n1331), .C2(n3212), .A(n4113), 
        .ZN(n4112) );
  AOI22_X1 U1841 ( .A1(n3165), .A2(n[1670]), .B1(n3160), .B2(n[1678]), .ZN(
        n4114) );
  OAI21_X1 U1842 ( .B1(n4131), .B2(n4132), .A(n3698), .ZN(n4130) );
  OAI221_X1 U1843 ( .B1(n1403), .B2(n3187), .C1(n1395), .C2(n3174), .A(n4134), 
        .ZN(n4131) );
  OAI221_X1 U1844 ( .B1(n1467), .B2(n3222), .C1(n1459), .C2(n3215), .A(n4133), 
        .ZN(n4132) );
  AOI22_X1 U1845 ( .A1(n3165), .A2(n[1606]), .B1(n3161), .B2(n[1614]), .ZN(
        n4134) );
  OAI21_X1 U1846 ( .B1(n4153), .B2(n4154), .A(n3666), .ZN(n4152) );
  OAI221_X1 U1847 ( .B1(n411), .B2(n3186), .C1(n403), .C2(n3173), .A(n4156), 
        .ZN(n4153) );
  OAI221_X1 U1848 ( .B1(n443), .B2(n3221), .C1(n435), .C2(n3209), .A(n4155), 
        .ZN(n4154) );
  AOI22_X1 U1849 ( .A1(n3164), .A2(n[2182]), .B1(n3161), .B2(n[2190]), .ZN(
        n4156) );
  OAI21_X1 U1850 ( .B1(n4173), .B2(n4174), .A(n3698), .ZN(n4172) );
  OAI221_X1 U1851 ( .B1(n475), .B2(n3186), .C1(n467), .C2(n3178), .A(n4176), 
        .ZN(n4173) );
  OAI221_X1 U1852 ( .B1(n507), .B2(n3221), .C1(n499), .C2(n3214), .A(n4175), 
        .ZN(n4174) );
  AOI22_X1 U1853 ( .A1(n3164), .A2(n[2118]), .B1(n3156), .B2(n[2126]), .ZN(
        n4176) );
  OAI21_X1 U1854 ( .B1(n3959), .B2(n3960), .A(n3698), .ZN(n3958) );
  OAI221_X1 U1855 ( .B1(n1402), .B2(n3189), .C1(n1394), .C2(n3175), .A(n3962), 
        .ZN(n3959) );
  OAI221_X1 U1856 ( .B1(n1466), .B2(n3224), .C1(n1458), .C2(n3212), .A(n3961), 
        .ZN(n3960) );
  AOI22_X1 U1857 ( .A1(n3167), .A2(n[1607]), .B1(n3156), .B2(n[1615]), .ZN(
        n3962) );
  OAI21_X1 U1858 ( .B1(n3981), .B2(n3982), .A(n3666), .ZN(n3980) );
  OAI221_X1 U1859 ( .B1(n410), .B2(n3189), .C1(n402), .C2(n3175), .A(n3984), 
        .ZN(n3981) );
  OAI221_X1 U1860 ( .B1(n442), .B2(n3224), .C1(n434), .C2(n3212), .A(n3983), 
        .ZN(n3982) );
  AOI22_X1 U1861 ( .A1(n3167), .A2(n[2183]), .B1(n3156), .B2(n[2191]), .ZN(
        n3984) );
  OAI21_X1 U1862 ( .B1(n4001), .B2(n4002), .A(n3698), .ZN(n4000) );
  OAI221_X1 U1863 ( .B1(n474), .B2(n3189), .C1(n466), .C2(n3175), .A(n4004), 
        .ZN(n4001) );
  OAI221_X1 U1864 ( .B1(n506), .B2(n3224), .C1(n498), .C2(n3212), .A(n4003), 
        .ZN(n4002) );
  AOI22_X1 U1865 ( .A1(n3167), .A2(n[2119]), .B1(n3156), .B2(n[2127]), .ZN(
        n4004) );
  OAI21_X1 U1866 ( .B1(n4891), .B2(n4892), .A(n3152), .ZN(n4885) );
  OAI221_X1 U1867 ( .B1(n2848), .B2(n3181), .C1(n2840), .C2(n3175), .A(n4894), 
        .ZN(n4891) );
  OAI221_X1 U1868 ( .B1(n2880), .B2(n3225), .C1(n2872), .C2(n3668), .A(n4893), 
        .ZN(n4892) );
  AOI22_X1 U1869 ( .A1(n3167), .A2(n[769]), .B1(n3676), .B2(n[777]), .ZN(n4894) );
  OAI21_X1 U1870 ( .B1(n4911), .B2(n4912), .A(n3703), .ZN(n4905) );
  OAI221_X1 U1871 ( .B1(n2912), .B2(n3189), .C1(n2904), .C2(n3673), .A(n4914), 
        .ZN(n4911) );
  OAI221_X1 U1872 ( .B1(n2944), .B2(n3223), .C1(n2936), .C2(n3668), .A(n4913), 
        .ZN(n4912) );
  AOI22_X1 U1873 ( .A1(n3170), .A2(n[705]), .B1(n3153), .B2(n[713]), .ZN(n4914) );
  OAI21_X1 U1874 ( .B1(n4719), .B2(n4720), .A(n3152), .ZN(n4713) );
  OAI221_X1 U1875 ( .B1(n2847), .B2(n3181), .C1(n2839), .C2(n3673), .A(n4722), 
        .ZN(n4719) );
  OAI221_X1 U1876 ( .B1(n2879), .B2(n3218), .C1(n2871), .C2(n3214), .A(n4721), 
        .ZN(n4720) );
  AOI22_X1 U1877 ( .A1(n3164), .A2(n[770]), .B1(n3155), .B2(n[778]), .ZN(n4722) );
  OAI21_X1 U1878 ( .B1(n4739), .B2(n4740), .A(n3703), .ZN(n4733) );
  OAI221_X1 U1879 ( .B1(n2911), .B2(n3184), .C1(n2903), .C2(n3180), .A(n4742), 
        .ZN(n4739) );
  OAI221_X1 U1880 ( .B1(n2943), .B2(n3223), .C1(n2935), .C2(n3209), .A(n4741), 
        .ZN(n4740) );
  AOI22_X1 U1881 ( .A1(n3167), .A2(n[706]), .B1(n3153), .B2(n[714]), .ZN(n4742) );
  OAI21_X1 U1882 ( .B1(n4203), .B2(n4204), .A(n3679), .ZN(n4197) );
  OAI221_X1 U1883 ( .B1(n2844), .B2(n3186), .C1(n2836), .C2(n3178), .A(n4206), 
        .ZN(n4203) );
  OAI221_X1 U1884 ( .B1(n2876), .B2(n3221), .C1(n2868), .C2(n3215), .A(n4205), 
        .ZN(n4204) );
  AOI22_X1 U1885 ( .A1(n3164), .A2(n[773]), .B1(n3155), .B2(n[781]), .ZN(n4206) );
  OAI21_X1 U1886 ( .B1(n4223), .B2(n4224), .A(n3148), .ZN(n4217) );
  OAI221_X1 U1887 ( .B1(n2908), .B2(n3185), .C1(n2900), .C2(n3174), .A(n4226), 
        .ZN(n4223) );
  OAI221_X1 U1888 ( .B1(n2940), .B2(n3220), .C1(n2932), .C2(n3211), .A(n4225), 
        .ZN(n4224) );
  AOI22_X1 U1889 ( .A1(n3163), .A2(n[709]), .B1(n3155), .B2(n[717]), .ZN(n4226) );
  OAI21_X1 U1890 ( .B1(n4031), .B2(n4032), .A(n3152), .ZN(n4025) );
  OAI221_X1 U1891 ( .B1(n2843), .B2(n3188), .C1(n2835), .C2(n3177), .A(n4034), 
        .ZN(n4031) );
  OAI221_X1 U1892 ( .B1(n2875), .B2(n3223), .C1(n2867), .C2(n3216), .A(n4033), 
        .ZN(n4032) );
  AOI22_X1 U1893 ( .A1(n3166), .A2(n[774]), .B1(n3158), .B2(n[782]), .ZN(n4034) );
  OAI21_X1 U1894 ( .B1(n4051), .B2(n4052), .A(n3703), .ZN(n4045) );
  OAI221_X1 U1895 ( .B1(n2907), .B2(n3188), .C1(n2899), .C2(n3177), .A(n4054), 
        .ZN(n4051) );
  OAI221_X1 U1896 ( .B1(n2939), .B2(n3223), .C1(n2931), .C2(n3212), .A(n4053), 
        .ZN(n4052) );
  AOI22_X1 U1897 ( .A1(n3166), .A2(n[710]), .B1(n3158), .B2(n[718]), .ZN(n4054) );
  OAI22_X1 U1898 ( .A1(n3145), .A2(n3652), .B1(n3297), .B2(n1984), .ZN(n5824)
         );
  OAI22_X1 U1899 ( .A1(n3132), .A2(n3652), .B1(n3297), .B2(n1983), .ZN(n5825)
         );
  OAI22_X1 U1900 ( .A1(n3119), .A2(n3652), .B1(n3297), .B2(n1982), .ZN(n5826)
         );
  OAI22_X1 U1901 ( .A1(n3117), .A2(n3652), .B1(n3297), .B2(n1981), .ZN(n5827)
         );
  OAI22_X1 U1902 ( .A1(n3104), .A2(n3652), .B1(n3297), .B2(n1980), .ZN(n5828)
         );
  OAI22_X1 U1903 ( .A1(n3094), .A2(n3652), .B1(n3297), .B2(n1979), .ZN(n5829)
         );
  OAI22_X1 U1904 ( .A1(n3090), .A2(n3652), .B1(n3297), .B2(n1978), .ZN(n5830)
         );
  OAI22_X1 U1905 ( .A1(n3081), .A2(n3652), .B1(n3297), .B2(n1977), .ZN(n5831)
         );
  OAI22_X1 U1906 ( .A1(n3140), .A2(n3353), .B1(n7244), .B2(n1944), .ZN(n5848)
         );
  OAI22_X1 U1907 ( .A1(n7257), .A2(n3353), .B1(n7244), .B2(n1943), .ZN(n5849)
         );
  OAI22_X1 U1908 ( .A1(n3121), .A2(n3353), .B1(n7244), .B2(n1942), .ZN(n5850)
         );
  OAI22_X1 U1909 ( .A1(n7255), .A2(n3353), .B1(n7244), .B2(n1941), .ZN(n5851)
         );
  OAI22_X1 U1910 ( .A1(n3106), .A2(n3353), .B1(n7244), .B2(n1940), .ZN(n5852)
         );
  OAI22_X1 U1911 ( .A1(n3091), .A2(n3353), .B1(n7244), .B2(n1939), .ZN(n5853)
         );
  OAI22_X1 U1912 ( .A1(n3084), .A2(n3353), .B1(n7244), .B2(n1938), .ZN(n5854)
         );
  OAI22_X1 U1913 ( .A1(n3075), .A2(n3353), .B1(n7244), .B2(n1937), .ZN(n5855)
         );
  OAI22_X1 U1914 ( .A1(n3139), .A2(n3355), .B1(n7115), .B2(n1920), .ZN(n5856)
         );
  OAI22_X1 U1915 ( .A1(n7257), .A2(n3355), .B1(n7115), .B2(n1919), .ZN(n5857)
         );
  OAI22_X1 U1916 ( .A1(n3121), .A2(n3355), .B1(n7115), .B2(n1918), .ZN(n5858)
         );
  OAI22_X1 U1917 ( .A1(n3109), .A2(n3355), .B1(n7115), .B2(n1917), .ZN(n5859)
         );
  OAI22_X1 U1918 ( .A1(n7254), .A2(n3355), .B1(n7115), .B2(n1916), .ZN(n5860)
         );
  OAI22_X1 U1919 ( .A1(n7253), .A2(n3355), .B1(n7115), .B2(n1915), .ZN(n5861)
         );
  OAI22_X1 U1920 ( .A1(n3087), .A2(n3355), .B1(n7115), .B2(n1914), .ZN(n5862)
         );
  OAI22_X1 U1921 ( .A1(n3078), .A2(n3355), .B1(n7115), .B2(n1913), .ZN(n5863)
         );
  OAI22_X1 U1922 ( .A1(n3140), .A2(n3357), .B1(n7180), .B2(n1912), .ZN(n5864)
         );
  OAI22_X1 U1923 ( .A1(n7257), .A2(n3357), .B1(n7180), .B2(n1911), .ZN(n5865)
         );
  OAI22_X1 U1924 ( .A1(n3121), .A2(n3357), .B1(n7180), .B2(n1910), .ZN(n5866)
         );
  OAI22_X1 U1925 ( .A1(n3109), .A2(n3357), .B1(n7180), .B2(n1909), .ZN(n5867)
         );
  OAI22_X1 U1926 ( .A1(n7254), .A2(n3357), .B1(n7180), .B2(n1908), .ZN(n5868)
         );
  OAI22_X1 U1927 ( .A1(n3096), .A2(n3357), .B1(n7180), .B2(n1907), .ZN(n5869)
         );
  OAI22_X1 U1928 ( .A1(n3089), .A2(n3357), .B1(n7180), .B2(n1906), .ZN(n5870)
         );
  OAI22_X1 U1929 ( .A1(n3080), .A2(n3357), .B1(n7180), .B2(n1905), .ZN(n5871)
         );
  OAI22_X1 U1930 ( .A1(n3139), .A2(n3359), .B1(n3280), .B2(n1888), .ZN(n5872)
         );
  OAI22_X1 U1931 ( .A1(n7257), .A2(n3359), .B1(n3280), .B2(n1887), .ZN(n5873)
         );
  OAI22_X1 U1932 ( .A1(n3121), .A2(n3359), .B1(n3280), .B2(n1886), .ZN(n5874)
         );
  OAI22_X1 U1933 ( .A1(n3117), .A2(n3359), .B1(n3280), .B2(n1885), .ZN(n5875)
         );
  OAI22_X1 U1934 ( .A1(n7254), .A2(n3359), .B1(n3280), .B2(n1884), .ZN(n5876)
         );
  OAI22_X1 U1935 ( .A1(n3091), .A2(n3359), .B1(n3280), .B2(n1883), .ZN(n5877)
         );
  OAI22_X1 U1936 ( .A1(n3085), .A2(n3359), .B1(n3280), .B2(n1882), .ZN(n5878)
         );
  OAI22_X1 U1937 ( .A1(n3076), .A2(n3359), .B1(n3280), .B2(n1881), .ZN(n5879)
         );
  OAI22_X1 U1938 ( .A1(n3140), .A2(n3361), .B1(n7228), .B2(n1880), .ZN(n5880)
         );
  OAI22_X1 U1939 ( .A1(n7257), .A2(n3361), .B1(n7228), .B2(n1879), .ZN(n5881)
         );
  OAI22_X1 U1940 ( .A1(n3121), .A2(n3361), .B1(n7228), .B2(n1878), .ZN(n5882)
         );
  OAI22_X1 U1941 ( .A1(n7255), .A2(n3361), .B1(n7228), .B2(n1877), .ZN(n5883)
         );
  OAI22_X1 U1942 ( .A1(n7254), .A2(n3361), .B1(n7228), .B2(n1876), .ZN(n5884)
         );
  OAI22_X1 U1943 ( .A1(n3096), .A2(n3361), .B1(n7228), .B2(n1875), .ZN(n5885)
         );
  OAI22_X1 U1944 ( .A1(n7252), .A2(n3361), .B1(n7228), .B2(n1874), .ZN(n5886)
         );
  OAI22_X1 U1945 ( .A1(n7251), .A2(n3361), .B1(n7228), .B2(n1873), .ZN(n5887)
         );
  OAI22_X1 U1946 ( .A1(n3139), .A2(n3363), .B1(n3344), .B2(n1856), .ZN(n5888)
         );
  OAI22_X1 U1947 ( .A1(n7257), .A2(n3363), .B1(n3344), .B2(n1855), .ZN(n5889)
         );
  OAI22_X1 U1948 ( .A1(n3121), .A2(n3363), .B1(n3344), .B2(n1854), .ZN(n5890)
         );
  OAI22_X1 U1949 ( .A1(n7255), .A2(n3363), .B1(n3344), .B2(n1853), .ZN(n5891)
         );
  OAI22_X1 U1950 ( .A1(n7254), .A2(n3363), .B1(n3344), .B2(n1852), .ZN(n5892)
         );
  OAI22_X1 U1951 ( .A1(n3091), .A2(n3363), .B1(n3344), .B2(n1851), .ZN(n5893)
         );
  OAI22_X1 U1952 ( .A1(n7252), .A2(n3363), .B1(n3344), .B2(n1850), .ZN(n5894)
         );
  OAI22_X1 U1953 ( .A1(n7251), .A2(n3363), .B1(n3344), .B2(n1849), .ZN(n5895)
         );
  OAI22_X1 U1954 ( .A1(n3140), .A2(n3365), .B1(n7164), .B2(n1848), .ZN(n5896)
         );
  OAI22_X1 U1955 ( .A1(n7257), .A2(n3365), .B1(n7164), .B2(n1847), .ZN(n5897)
         );
  OAI22_X1 U1956 ( .A1(n3121), .A2(n3365), .B1(n7164), .B2(n1846), .ZN(n5898)
         );
  OAI22_X1 U1957 ( .A1(n7255), .A2(n3365), .B1(n7164), .B2(n1845), .ZN(n5899)
         );
  OAI22_X1 U1958 ( .A1(n7254), .A2(n3365), .B1(n7164), .B2(n1844), .ZN(n5900)
         );
  OAI22_X1 U1959 ( .A1(n3098), .A2(n3365), .B1(n7164), .B2(n1843), .ZN(n5901)
         );
  OAI22_X1 U1960 ( .A1(n7252), .A2(n3365), .B1(n7164), .B2(n1842), .ZN(n5902)
         );
  OAI22_X1 U1961 ( .A1(n7251), .A2(n3365), .B1(n7164), .B2(n1841), .ZN(n5903)
         );
  OAI22_X1 U1962 ( .A1(n3139), .A2(n3367), .B1(n3264), .B2(n1824), .ZN(n5904)
         );
  OAI22_X1 U1963 ( .A1(n7257), .A2(n3367), .B1(n3264), .B2(n1823), .ZN(n5905)
         );
  OAI22_X1 U1964 ( .A1(n3121), .A2(n3367), .B1(n3264), .B2(n1822), .ZN(n5906)
         );
  OAI22_X1 U1965 ( .A1(n7255), .A2(n3367), .B1(n3264), .B2(n1821), .ZN(n5907)
         );
  OAI22_X1 U1966 ( .A1(n7254), .A2(n3367), .B1(n3264), .B2(n1820), .ZN(n5908)
         );
  OAI22_X1 U1967 ( .A1(n3091), .A2(n3367), .B1(n3264), .B2(n1819), .ZN(n5909)
         );
  OAI22_X1 U1968 ( .A1(n7252), .A2(n3367), .B1(n3264), .B2(n1818), .ZN(n5910)
         );
  OAI22_X1 U1969 ( .A1(n7251), .A2(n3367), .B1(n3264), .B2(n1817), .ZN(n5911)
         );
  OAI22_X1 U1970 ( .A1(n3140), .A2(n3369), .B1(n7212), .B2(n1816), .ZN(n5912)
         );
  OAI22_X1 U1971 ( .A1(n7257), .A2(n3369), .B1(n7212), .B2(n1815), .ZN(n5913)
         );
  OAI22_X1 U1972 ( .A1(n3121), .A2(n3369), .B1(n7212), .B2(n1814), .ZN(n5914)
         );
  OAI22_X1 U1973 ( .A1(n7255), .A2(n3369), .B1(n7212), .B2(n1813), .ZN(n5915)
         );
  OAI22_X1 U1974 ( .A1(n7254), .A2(n3369), .B1(n7212), .B2(n1812), .ZN(n5916)
         );
  OAI22_X1 U1975 ( .A1(n3099), .A2(n3369), .B1(n7212), .B2(n1811), .ZN(n5917)
         );
  OAI22_X1 U1976 ( .A1(n7252), .A2(n3369), .B1(n7212), .B2(n1810), .ZN(n5918)
         );
  OAI22_X1 U1977 ( .A1(n7251), .A2(n3369), .B1(n7212), .B2(n1809), .ZN(n5919)
         );
  OAI22_X1 U1978 ( .A1(n3139), .A2(n3371), .B1(n3328), .B2(n1792), .ZN(n5920)
         );
  OAI22_X1 U1979 ( .A1(n3131), .A2(n3371), .B1(n3328), .B2(n1791), .ZN(n5921)
         );
  OAI22_X1 U1980 ( .A1(n3120), .A2(n3371), .B1(n3328), .B2(n1790), .ZN(n5922)
         );
  OAI22_X1 U1981 ( .A1(n7255), .A2(n3371), .B1(n3328), .B2(n1789), .ZN(n5923)
         );
  OAI22_X1 U1982 ( .A1(n7254), .A2(n3371), .B1(n3328), .B2(n1788), .ZN(n5924)
         );
  OAI22_X1 U1983 ( .A1(n3091), .A2(n3371), .B1(n3328), .B2(n1787), .ZN(n5925)
         );
  OAI22_X1 U1984 ( .A1(n7252), .A2(n3371), .B1(n3328), .B2(n1786), .ZN(n5926)
         );
  OAI22_X1 U1985 ( .A1(n7251), .A2(n3371), .B1(n3328), .B2(n1785), .ZN(n5927)
         );
  OAI22_X1 U1986 ( .A1(n3140), .A2(n3373), .B1(n7148), .B2(n1784), .ZN(n5928)
         );
  OAI22_X1 U1987 ( .A1(n3129), .A2(n3373), .B1(n7148), .B2(n1783), .ZN(n5929)
         );
  OAI22_X1 U1988 ( .A1(n3121), .A2(n3373), .B1(n7148), .B2(n1782), .ZN(n5930)
         );
  OAI22_X1 U1989 ( .A1(n7255), .A2(n3373), .B1(n7148), .B2(n1781), .ZN(n5931)
         );
  OAI22_X1 U1990 ( .A1(n7254), .A2(n3373), .B1(n7148), .B2(n1780), .ZN(n5932)
         );
  OAI22_X1 U1991 ( .A1(n3097), .A2(n3373), .B1(n7148), .B2(n1779), .ZN(n5933)
         );
  OAI22_X1 U1992 ( .A1(n7252), .A2(n3373), .B1(n7148), .B2(n1778), .ZN(n5934)
         );
  OAI22_X1 U1993 ( .A1(n7251), .A2(n3373), .B1(n7148), .B2(n1777), .ZN(n5935)
         );
  OAI22_X1 U1994 ( .A1(n7258), .A2(n3375), .B1(n3248), .B2(n1760), .ZN(n5936)
         );
  OAI22_X1 U1995 ( .A1(n3130), .A2(n3375), .B1(n3248), .B2(n1759), .ZN(n5937)
         );
  OAI22_X1 U1996 ( .A1(n3120), .A2(n3375), .B1(n3248), .B2(n1758), .ZN(n5938)
         );
  OAI22_X1 U1997 ( .A1(n3117), .A2(n3375), .B1(n3248), .B2(n1757), .ZN(n5939)
         );
  OAI22_X1 U1998 ( .A1(n7254), .A2(n3375), .B1(n3248), .B2(n1756), .ZN(n5940)
         );
  OAI22_X1 U1999 ( .A1(n3098), .A2(n3375), .B1(n3248), .B2(n1755), .ZN(n5941)
         );
  OAI22_X1 U2000 ( .A1(n3085), .A2(n3375), .B1(n3248), .B2(n1754), .ZN(n5942)
         );
  OAI22_X1 U2001 ( .A1(n3076), .A2(n3375), .B1(n3248), .B2(n1753), .ZN(n5943)
         );
  OAI22_X1 U2002 ( .A1(n3145), .A2(n3377), .B1(n7196), .B2(n1752), .ZN(n5944)
         );
  OAI22_X1 U2003 ( .A1(n3129), .A2(n3377), .B1(n7196), .B2(n1751), .ZN(n5945)
         );
  OAI22_X1 U2004 ( .A1(n3119), .A2(n3377), .B1(n7196), .B2(n1750), .ZN(n5946)
         );
  OAI22_X1 U2005 ( .A1(n3116), .A2(n3377), .B1(n7196), .B2(n1749), .ZN(n5947)
         );
  OAI22_X1 U2006 ( .A1(n3106), .A2(n3377), .B1(n7196), .B2(n1748), .ZN(n5948)
         );
  OAI22_X1 U2007 ( .A1(n3093), .A2(n3377), .B1(n7196), .B2(n1747), .ZN(n5949)
         );
  OAI22_X1 U2008 ( .A1(n3084), .A2(n3377), .B1(n7196), .B2(n1746), .ZN(n5950)
         );
  OAI22_X1 U2009 ( .A1(n3075), .A2(n3377), .B1(n7196), .B2(n1745), .ZN(n5951)
         );
  OAI22_X1 U2010 ( .A1(n3138), .A2(n3379), .B1(n3312), .B2(n1728), .ZN(n5952)
         );
  OAI22_X1 U2011 ( .A1(n3129), .A2(n3379), .B1(n3312), .B2(n1727), .ZN(n5953)
         );
  OAI22_X1 U2012 ( .A1(n3119), .A2(n3379), .B1(n3312), .B2(n1726), .ZN(n5954)
         );
  OAI22_X1 U2013 ( .A1(n3117), .A2(n3379), .B1(n3312), .B2(n1725), .ZN(n5955)
         );
  OAI22_X1 U2014 ( .A1(n3106), .A2(n3379), .B1(n3312), .B2(n1724), .ZN(n5956)
         );
  OAI22_X1 U2015 ( .A1(n3098), .A2(n3379), .B1(n3312), .B2(n1723), .ZN(n5957)
         );
  OAI22_X1 U2016 ( .A1(n3090), .A2(n3379), .B1(n3312), .B2(n1722), .ZN(n5958)
         );
  OAI22_X1 U2017 ( .A1(n3081), .A2(n3379), .B1(n3312), .B2(n1721), .ZN(n5959)
         );
  OAI22_X1 U2018 ( .A1(n3143), .A2(n3541), .B1(n3303), .B2(n3072), .ZN(n5056)
         );
  OAI22_X1 U2019 ( .A1(n3135), .A2(n3541), .B1(n3303), .B2(n3071), .ZN(n5057)
         );
  OAI22_X1 U2020 ( .A1(n3125), .A2(n3541), .B1(n3303), .B2(n3070), .ZN(n5058)
         );
  OAI22_X1 U2021 ( .A1(n3112), .A2(n3541), .B1(n3303), .B2(n3069), .ZN(n5059)
         );
  OAI22_X1 U2022 ( .A1(n3102), .A2(n3541), .B1(n3303), .B2(n3068), .ZN(n5060)
         );
  OAI22_X1 U2023 ( .A1(n3096), .A2(n3541), .B1(n3303), .B2(n3067), .ZN(n5061)
         );
  OAI22_X1 U2024 ( .A1(n3087), .A2(n3541), .B1(n3303), .B2(n3066), .ZN(n5062)
         );
  OAI22_X1 U2025 ( .A1(n3078), .A2(n3541), .B1(n3303), .B2(n3065), .ZN(n5063)
         );
  OAI22_X1 U2026 ( .A1(n3143), .A2(n3543), .B1(n7123), .B2(n3064), .ZN(n5064)
         );
  OAI22_X1 U2027 ( .A1(n3135), .A2(n3543), .B1(n7123), .B2(n3063), .ZN(n5065)
         );
  OAI22_X1 U2028 ( .A1(n3125), .A2(n3543), .B1(n7123), .B2(n3062), .ZN(n5066)
         );
  OAI22_X1 U2029 ( .A1(n3113), .A2(n3543), .B1(n7123), .B2(n3061), .ZN(n5067)
         );
  OAI22_X1 U2030 ( .A1(n3102), .A2(n3543), .B1(n7123), .B2(n3060), .ZN(n5068)
         );
  OAI22_X1 U2031 ( .A1(n3096), .A2(n3543), .B1(n7123), .B2(n3059), .ZN(n5069)
         );
  OAI22_X1 U2032 ( .A1(n3087), .A2(n3543), .B1(n7123), .B2(n3058), .ZN(n5070)
         );
  OAI22_X1 U2033 ( .A1(n3078), .A2(n3543), .B1(n7123), .B2(n3057), .ZN(n5071)
         );
  OAI22_X1 U2034 ( .A1(n3143), .A2(n3544), .B1(n3286), .B2(n3056), .ZN(n5072)
         );
  OAI22_X1 U2035 ( .A1(n3135), .A2(n3544), .B1(n3286), .B2(n3055), .ZN(n5073)
         );
  OAI22_X1 U2036 ( .A1(n3125), .A2(n3544), .B1(n3286), .B2(n3054), .ZN(n5074)
         );
  OAI22_X1 U2037 ( .A1(n3114), .A2(n3544), .B1(n3286), .B2(n3053), .ZN(n5075)
         );
  OAI22_X1 U2038 ( .A1(n3102), .A2(n3544), .B1(n3286), .B2(n3052), .ZN(n5076)
         );
  OAI22_X1 U2039 ( .A1(n3096), .A2(n3544), .B1(n3286), .B2(n3051), .ZN(n5077)
         );
  OAI22_X1 U2040 ( .A1(n3087), .A2(n3544), .B1(n3286), .B2(n3050), .ZN(n5078)
         );
  OAI22_X1 U2041 ( .A1(n3078), .A2(n3544), .B1(n3286), .B2(n3049), .ZN(n5079)
         );
  OAI22_X1 U2042 ( .A1(n3143), .A2(n3545), .B1(n7234), .B2(n3048), .ZN(n5080)
         );
  OAI22_X1 U2043 ( .A1(n3135), .A2(n3545), .B1(n7234), .B2(n3047), .ZN(n5081)
         );
  OAI22_X1 U2044 ( .A1(n3125), .A2(n3545), .B1(n7234), .B2(n3046), .ZN(n5082)
         );
  OAI22_X1 U2045 ( .A1(n3115), .A2(n3545), .B1(n7234), .B2(n3045), .ZN(n5083)
         );
  OAI22_X1 U2046 ( .A1(n3102), .A2(n3545), .B1(n7234), .B2(n3044), .ZN(n5084)
         );
  OAI22_X1 U2047 ( .A1(n3096), .A2(n3545), .B1(n7234), .B2(n3043), .ZN(n5085)
         );
  OAI22_X1 U2048 ( .A1(n3087), .A2(n3545), .B1(n7234), .B2(n3042), .ZN(n5086)
         );
  OAI22_X1 U2049 ( .A1(n3078), .A2(n3545), .B1(n7234), .B2(n3041), .ZN(n5087)
         );
  OAI22_X1 U2050 ( .A1(n3142), .A2(n3546), .B1(n7105), .B2(n3040), .ZN(n5088)
         );
  OAI22_X1 U2051 ( .A1(n3133), .A2(n3546), .B1(n7105), .B2(n3039), .ZN(n5089)
         );
  OAI22_X1 U2052 ( .A1(n3124), .A2(n3546), .B1(n7105), .B2(n3038), .ZN(n5090)
         );
  OAI22_X1 U2053 ( .A1(n3112), .A2(n3546), .B1(n7105), .B2(n3037), .ZN(n5091)
         );
  OAI22_X1 U2054 ( .A1(n3102), .A2(n3546), .B1(n7105), .B2(n3036), .ZN(n5092)
         );
  OAI22_X1 U2055 ( .A1(n3096), .A2(n3546), .B1(n7105), .B2(n3035), .ZN(n5093)
         );
  OAI22_X1 U2056 ( .A1(n3087), .A2(n3546), .B1(n7105), .B2(n3034), .ZN(n5094)
         );
  OAI22_X1 U2057 ( .A1(n3078), .A2(n3546), .B1(n7105), .B2(n3033), .ZN(n5095)
         );
  OAI22_X1 U2058 ( .A1(n3142), .A2(n3547), .B1(n7170), .B2(n3032), .ZN(n5096)
         );
  OAI22_X1 U2059 ( .A1(n3135), .A2(n3547), .B1(n7170), .B2(n3031), .ZN(n5097)
         );
  OAI22_X1 U2060 ( .A1(n3124), .A2(n3547), .B1(n7170), .B2(n3030), .ZN(n5098)
         );
  OAI22_X1 U2061 ( .A1(n3113), .A2(n3547), .B1(n7170), .B2(n3029), .ZN(n5099)
         );
  OAI22_X1 U2062 ( .A1(n3102), .A2(n3547), .B1(n7170), .B2(n3028), .ZN(n5100)
         );
  OAI22_X1 U2063 ( .A1(n3096), .A2(n3547), .B1(n7170), .B2(n3027), .ZN(n5101)
         );
  OAI22_X1 U2064 ( .A1(n3087), .A2(n3547), .B1(n7170), .B2(n3026), .ZN(n5102)
         );
  OAI22_X1 U2065 ( .A1(n3078), .A2(n3547), .B1(n7170), .B2(n3025), .ZN(n5103)
         );
  OAI22_X1 U2066 ( .A1(n3142), .A2(n3548), .B1(n3270), .B2(n3024), .ZN(n5104)
         );
  OAI22_X1 U2067 ( .A1(n3136), .A2(n3548), .B1(n3270), .B2(n3023), .ZN(n5105)
         );
  OAI22_X1 U2068 ( .A1(n3124), .A2(n3548), .B1(n3270), .B2(n3022), .ZN(n5106)
         );
  OAI22_X1 U2069 ( .A1(n3114), .A2(n3548), .B1(n3270), .B2(n3021), .ZN(n5107)
         );
  OAI22_X1 U2070 ( .A1(n3102), .A2(n3548), .B1(n3270), .B2(n3020), .ZN(n5108)
         );
  OAI22_X1 U2071 ( .A1(n3096), .A2(n3548), .B1(n3270), .B2(n3019), .ZN(n5109)
         );
  OAI22_X1 U2072 ( .A1(n3087), .A2(n3548), .B1(n3270), .B2(n3018), .ZN(n5110)
         );
  OAI22_X1 U2073 ( .A1(n3078), .A2(n3548), .B1(n3270), .B2(n3017), .ZN(n5111)
         );
  OAI22_X1 U2074 ( .A1(n3142), .A2(n3549), .B1(n7218), .B2(n3016), .ZN(n5112)
         );
  OAI22_X1 U2075 ( .A1(n3132), .A2(n3549), .B1(n7218), .B2(n3015), .ZN(n5113)
         );
  OAI22_X1 U2076 ( .A1(n3124), .A2(n3549), .B1(n7218), .B2(n3014), .ZN(n5114)
         );
  OAI22_X1 U2077 ( .A1(n3115), .A2(n3549), .B1(n7218), .B2(n3013), .ZN(n5115)
         );
  OAI22_X1 U2078 ( .A1(n3102), .A2(n3549), .B1(n7218), .B2(n3012), .ZN(n5116)
         );
  OAI22_X1 U2079 ( .A1(n3096), .A2(n3549), .B1(n7218), .B2(n3011), .ZN(n5117)
         );
  OAI22_X1 U2080 ( .A1(n3087), .A2(n3549), .B1(n7218), .B2(n3010), .ZN(n5118)
         );
  OAI22_X1 U2081 ( .A1(n3078), .A2(n3549), .B1(n7218), .B2(n3009), .ZN(n5119)
         );
  OAI22_X1 U2082 ( .A1(n3142), .A2(n3550), .B1(n3334), .B2(n3008), .ZN(n5120)
         );
  OAI22_X1 U2083 ( .A1(n3131), .A2(n3550), .B1(n3334), .B2(n3007), .ZN(n5121)
         );
  OAI22_X1 U2084 ( .A1(n3124), .A2(n3550), .B1(n3334), .B2(n3006), .ZN(n5122)
         );
  OAI22_X1 U2085 ( .A1(n3112), .A2(n3550), .B1(n3334), .B2(n3005), .ZN(n5123)
         );
  OAI22_X1 U2086 ( .A1(n3102), .A2(n3550), .B1(n3334), .B2(n3004), .ZN(n5124)
         );
  OAI22_X1 U2087 ( .A1(n3096), .A2(n3550), .B1(n3334), .B2(n3003), .ZN(n5125)
         );
  OAI22_X1 U2088 ( .A1(n3087), .A2(n3550), .B1(n3334), .B2(n3002), .ZN(n5126)
         );
  OAI22_X1 U2089 ( .A1(n3078), .A2(n3550), .B1(n3334), .B2(n3001), .ZN(n5127)
         );
  OAI22_X1 U2090 ( .A1(n3142), .A2(n3551), .B1(n7154), .B2(n3000), .ZN(n5128)
         );
  OAI22_X1 U2091 ( .A1(n3134), .A2(n3551), .B1(n7154), .B2(n2999), .ZN(n5129)
         );
  OAI22_X1 U2092 ( .A1(n3124), .A2(n3551), .B1(n7154), .B2(n2998), .ZN(n5130)
         );
  OAI22_X1 U2093 ( .A1(n3113), .A2(n3551), .B1(n7154), .B2(n2997), .ZN(n5131)
         );
  OAI22_X1 U2094 ( .A1(n3102), .A2(n3551), .B1(n7154), .B2(n2996), .ZN(n5132)
         );
  OAI22_X1 U2095 ( .A1(n3096), .A2(n3551), .B1(n7154), .B2(n2995), .ZN(n5133)
         );
  OAI22_X1 U2096 ( .A1(n3087), .A2(n3551), .B1(n7154), .B2(n2994), .ZN(n5134)
         );
  OAI22_X1 U2097 ( .A1(n3078), .A2(n3551), .B1(n7154), .B2(n2993), .ZN(n5135)
         );
  OAI22_X1 U2098 ( .A1(n3142), .A2(n3552), .B1(n3254), .B2(n2992), .ZN(n5136)
         );
  OAI22_X1 U2099 ( .A1(n3134), .A2(n3552), .B1(n3254), .B2(n2991), .ZN(n5137)
         );
  OAI22_X1 U2100 ( .A1(n3124), .A2(n3552), .B1(n3254), .B2(n2990), .ZN(n5138)
         );
  OAI22_X1 U2101 ( .A1(n3114), .A2(n3552), .B1(n3254), .B2(n2989), .ZN(n5139)
         );
  OAI22_X1 U2102 ( .A1(n3103), .A2(n3552), .B1(n3254), .B2(n2988), .ZN(n5140)
         );
  OAI22_X1 U2103 ( .A1(n3097), .A2(n3552), .B1(n3254), .B2(n2987), .ZN(n5141)
         );
  OAI22_X1 U2104 ( .A1(n3088), .A2(n3552), .B1(n3254), .B2(n2986), .ZN(n5142)
         );
  OAI22_X1 U2105 ( .A1(n3079), .A2(n3552), .B1(n3254), .B2(n2985), .ZN(n5143)
         );
  OAI22_X1 U2106 ( .A1(n3142), .A2(n3553), .B1(n7202), .B2(n2984), .ZN(n5144)
         );
  OAI22_X1 U2107 ( .A1(n3133), .A2(n3553), .B1(n7202), .B2(n2983), .ZN(n5145)
         );
  OAI22_X1 U2108 ( .A1(n3124), .A2(n3553), .B1(n7202), .B2(n2982), .ZN(n5146)
         );
  OAI22_X1 U2109 ( .A1(n3114), .A2(n3553), .B1(n7202), .B2(n2981), .ZN(n5147)
         );
  OAI22_X1 U2110 ( .A1(n3103), .A2(n3553), .B1(n7202), .B2(n2980), .ZN(n5148)
         );
  OAI22_X1 U2111 ( .A1(n3094), .A2(n3553), .B1(n7202), .B2(n2979), .ZN(n5149)
         );
  OAI22_X1 U2112 ( .A1(n3088), .A2(n3553), .B1(n7202), .B2(n2978), .ZN(n5150)
         );
  OAI22_X1 U2113 ( .A1(n3079), .A2(n3553), .B1(n7202), .B2(n2977), .ZN(n5151)
         );
  OAI22_X1 U2114 ( .A1(n3142), .A2(n3554), .B1(n3318), .B2(n2976), .ZN(n5152)
         );
  OAI22_X1 U2115 ( .A1(n3135), .A2(n3554), .B1(n3318), .B2(n2975), .ZN(n5153)
         );
  OAI22_X1 U2116 ( .A1(n3124), .A2(n3554), .B1(n3318), .B2(n2974), .ZN(n5154)
         );
  OAI22_X1 U2117 ( .A1(n3114), .A2(n3554), .B1(n3318), .B2(n2973), .ZN(n5155)
         );
  OAI22_X1 U2118 ( .A1(n3103), .A2(n3554), .B1(n3318), .B2(n2972), .ZN(n5156)
         );
  OAI22_X1 U2119 ( .A1(n3095), .A2(n3554), .B1(n3318), .B2(n2971), .ZN(n5157)
         );
  OAI22_X1 U2120 ( .A1(n3088), .A2(n3554), .B1(n3318), .B2(n2970), .ZN(n5158)
         );
  OAI22_X1 U2121 ( .A1(n3079), .A2(n3554), .B1(n3318), .B2(n2969), .ZN(n5159)
         );
  OAI22_X1 U2122 ( .A1(n3142), .A2(n3555), .B1(n7138), .B2(n2968), .ZN(n5160)
         );
  OAI22_X1 U2123 ( .A1(n3136), .A2(n3555), .B1(n7138), .B2(n2967), .ZN(n5161)
         );
  OAI22_X1 U2124 ( .A1(n3124), .A2(n3555), .B1(n7138), .B2(n2966), .ZN(n5162)
         );
  OAI22_X1 U2125 ( .A1(n3114), .A2(n3555), .B1(n7138), .B2(n2965), .ZN(n5163)
         );
  OAI22_X1 U2126 ( .A1(n3103), .A2(n3555), .B1(n7138), .B2(n2964), .ZN(n5164)
         );
  OAI22_X1 U2127 ( .A1(n3096), .A2(n3555), .B1(n7138), .B2(n2963), .ZN(n5165)
         );
  OAI22_X1 U2128 ( .A1(n3088), .A2(n3555), .B1(n7138), .B2(n2962), .ZN(n5166)
         );
  OAI22_X1 U2129 ( .A1(n3079), .A2(n3555), .B1(n7138), .B2(n2961), .ZN(n5167)
         );
  OAI22_X1 U2130 ( .A1(n3142), .A2(n3556), .B1(n3238), .B2(n2960), .ZN(n5168)
         );
  OAI22_X1 U2131 ( .A1(n3134), .A2(n3556), .B1(n3238), .B2(n2959), .ZN(n5169)
         );
  OAI22_X1 U2132 ( .A1(n3124), .A2(n3556), .B1(n3238), .B2(n2958), .ZN(n5170)
         );
  OAI22_X1 U2133 ( .A1(n3114), .A2(n3556), .B1(n3238), .B2(n2957), .ZN(n5171)
         );
  OAI22_X1 U2134 ( .A1(n3103), .A2(n3556), .B1(n3238), .B2(n2956), .ZN(n5172)
         );
  OAI22_X1 U2135 ( .A1(n3096), .A2(n3556), .B1(n3238), .B2(n2955), .ZN(n5173)
         );
  OAI22_X1 U2136 ( .A1(n3088), .A2(n3556), .B1(n3238), .B2(n2954), .ZN(n5174)
         );
  OAI22_X1 U2137 ( .A1(n3079), .A2(n3556), .B1(n3238), .B2(n2953), .ZN(n5175)
         );
  OAI22_X1 U2138 ( .A1(n3142), .A2(n3557), .B1(n7186), .B2(n2952), .ZN(n5176)
         );
  OAI22_X1 U2139 ( .A1(n3133), .A2(n3557), .B1(n7186), .B2(n2951), .ZN(n5177)
         );
  OAI22_X1 U2140 ( .A1(n3124), .A2(n3557), .B1(n7186), .B2(n2950), .ZN(n5178)
         );
  OAI22_X1 U2141 ( .A1(n3114), .A2(n3557), .B1(n7186), .B2(n2949), .ZN(n5179)
         );
  OAI22_X1 U2142 ( .A1(n3103), .A2(n3557), .B1(n7186), .B2(n2948), .ZN(n5180)
         );
  OAI22_X1 U2143 ( .A1(n3097), .A2(n3557), .B1(n7186), .B2(n2947), .ZN(n5181)
         );
  OAI22_X1 U2144 ( .A1(n3088), .A2(n3557), .B1(n7186), .B2(n2946), .ZN(n5182)
         );
  OAI22_X1 U2145 ( .A1(n3079), .A2(n3557), .B1(n7186), .B2(n2945), .ZN(n5183)
         );
  OAI22_X1 U2146 ( .A1(n3142), .A2(n3559), .B1(n3302), .B2(n2944), .ZN(n5184)
         );
  OAI22_X1 U2147 ( .A1(n3132), .A2(n3559), .B1(n3302), .B2(n2943), .ZN(n5185)
         );
  OAI22_X1 U2148 ( .A1(n3124), .A2(n3559), .B1(n3302), .B2(n2942), .ZN(n5186)
         );
  OAI22_X1 U2149 ( .A1(n3114), .A2(n3559), .B1(n3302), .B2(n2941), .ZN(n5187)
         );
  OAI22_X1 U2150 ( .A1(n3103), .A2(n3559), .B1(n3302), .B2(n2940), .ZN(n5188)
         );
  OAI22_X1 U2151 ( .A1(n3094), .A2(n3559), .B1(n3302), .B2(n2939), .ZN(n5189)
         );
  OAI22_X1 U2152 ( .A1(n3088), .A2(n3559), .B1(n3302), .B2(n2938), .ZN(n5190)
         );
  OAI22_X1 U2153 ( .A1(n3079), .A2(n3559), .B1(n3302), .B2(n2937), .ZN(n5191)
         );
  OAI22_X1 U2154 ( .A1(n3141), .A2(n3561), .B1(n7122), .B2(n2936), .ZN(n5192)
         );
  OAI22_X1 U2155 ( .A1(n3131), .A2(n3561), .B1(n7122), .B2(n2935), .ZN(n5193)
         );
  OAI22_X1 U2156 ( .A1(n3123), .A2(n3561), .B1(n7122), .B2(n2934), .ZN(n5194)
         );
  OAI22_X1 U2157 ( .A1(n3114), .A2(n3561), .B1(n7122), .B2(n2933), .ZN(n5195)
         );
  OAI22_X1 U2158 ( .A1(n3103), .A2(n3561), .B1(n7122), .B2(n2932), .ZN(n5196)
         );
  OAI22_X1 U2159 ( .A1(n3095), .A2(n3561), .B1(n7122), .B2(n2931), .ZN(n5197)
         );
  OAI22_X1 U2160 ( .A1(n3088), .A2(n3561), .B1(n7122), .B2(n2930), .ZN(n5198)
         );
  OAI22_X1 U2161 ( .A1(n3079), .A2(n3561), .B1(n7122), .B2(n2929), .ZN(n5199)
         );
  OAI22_X1 U2162 ( .A1(n3141), .A2(n3562), .B1(n3285), .B2(n2928), .ZN(n5200)
         );
  OAI22_X1 U2163 ( .A1(n3132), .A2(n3562), .B1(n3285), .B2(n2927), .ZN(n5201)
         );
  OAI22_X1 U2164 ( .A1(n3123), .A2(n3562), .B1(n3285), .B2(n2926), .ZN(n5202)
         );
  OAI22_X1 U2165 ( .A1(n3114), .A2(n3562), .B1(n3285), .B2(n2925), .ZN(n5203)
         );
  OAI22_X1 U2166 ( .A1(n3103), .A2(n3562), .B1(n3285), .B2(n2924), .ZN(n5204)
         );
  OAI22_X1 U2167 ( .A1(n3096), .A2(n3562), .B1(n3285), .B2(n2923), .ZN(n5205)
         );
  OAI22_X1 U2168 ( .A1(n3088), .A2(n3562), .B1(n3285), .B2(n2922), .ZN(n5206)
         );
  OAI22_X1 U2169 ( .A1(n3079), .A2(n3562), .B1(n3285), .B2(n2921), .ZN(n5207)
         );
  OAI22_X1 U2170 ( .A1(n3141), .A2(n3563), .B1(n7233), .B2(n2920), .ZN(n5208)
         );
  OAI22_X1 U2171 ( .A1(n3131), .A2(n3563), .B1(n7233), .B2(n2919), .ZN(n5209)
         );
  OAI22_X1 U2172 ( .A1(n3123), .A2(n3563), .B1(n7233), .B2(n2918), .ZN(n5210)
         );
  OAI22_X1 U2173 ( .A1(n3114), .A2(n3563), .B1(n7233), .B2(n2917), .ZN(n5211)
         );
  OAI22_X1 U2174 ( .A1(n3103), .A2(n3563), .B1(n7233), .B2(n2916), .ZN(n5212)
         );
  OAI22_X1 U2175 ( .A1(n3097), .A2(n3563), .B1(n7233), .B2(n2915), .ZN(n5213)
         );
  OAI22_X1 U2176 ( .A1(n3088), .A2(n3563), .B1(n7233), .B2(n2914), .ZN(n5214)
         );
  OAI22_X1 U2177 ( .A1(n3079), .A2(n3563), .B1(n7233), .B2(n2913), .ZN(n5215)
         );
  OAI22_X1 U2178 ( .A1(n3141), .A2(n3564), .B1(n7104), .B2(n2912), .ZN(n5216)
         );
  OAI22_X1 U2179 ( .A1(n3135), .A2(n3564), .B1(n7104), .B2(n2911), .ZN(n5217)
         );
  OAI22_X1 U2180 ( .A1(n3123), .A2(n3564), .B1(n7104), .B2(n2910), .ZN(n5218)
         );
  OAI22_X1 U2181 ( .A1(n3114), .A2(n3564), .B1(n7104), .B2(n2909), .ZN(n5219)
         );
  OAI22_X1 U2182 ( .A1(n3103), .A2(n3564), .B1(n7104), .B2(n2908), .ZN(n5220)
         );
  OAI22_X1 U2183 ( .A1(n3098), .A2(n3564), .B1(n7104), .B2(n2907), .ZN(n5221)
         );
  OAI22_X1 U2184 ( .A1(n3088), .A2(n3564), .B1(n7104), .B2(n2906), .ZN(n5222)
         );
  OAI22_X1 U2185 ( .A1(n3079), .A2(n3564), .B1(n7104), .B2(n2905), .ZN(n5223)
         );
  OAI22_X1 U2186 ( .A1(n3141), .A2(n3565), .B1(n7169), .B2(n2904), .ZN(n5224)
         );
  OAI22_X1 U2187 ( .A1(n3136), .A2(n3565), .B1(n7169), .B2(n2903), .ZN(n5225)
         );
  OAI22_X1 U2188 ( .A1(n3123), .A2(n3565), .B1(n7169), .B2(n2902), .ZN(n5226)
         );
  OAI22_X1 U2189 ( .A1(n3114), .A2(n3565), .B1(n7169), .B2(n2901), .ZN(n5227)
         );
  OAI22_X1 U2190 ( .A1(n3103), .A2(n3565), .B1(n7169), .B2(n2900), .ZN(n5228)
         );
  OAI22_X1 U2191 ( .A1(n3099), .A2(n3565), .B1(n7169), .B2(n2899), .ZN(n5229)
         );
  OAI22_X1 U2192 ( .A1(n3088), .A2(n3565), .B1(n7169), .B2(n2898), .ZN(n5230)
         );
  OAI22_X1 U2193 ( .A1(n3079), .A2(n3565), .B1(n7169), .B2(n2897), .ZN(n5231)
         );
  OAI22_X1 U2194 ( .A1(n3141), .A2(n3566), .B1(n3269), .B2(n2896), .ZN(n5232)
         );
  OAI22_X1 U2195 ( .A1(n3134), .A2(n3566), .B1(n3269), .B2(n2895), .ZN(n5233)
         );
  OAI22_X1 U2196 ( .A1(n3123), .A2(n3566), .B1(n3269), .B2(n2894), .ZN(n5234)
         );
  OAI22_X1 U2197 ( .A1(n3114), .A2(n3566), .B1(n3269), .B2(n2893), .ZN(n5235)
         );
  OAI22_X1 U2198 ( .A1(n3103), .A2(n3566), .B1(n3269), .B2(n2892), .ZN(n5236)
         );
  OAI22_X1 U2199 ( .A1(n3091), .A2(n3566), .B1(n3269), .B2(n2891), .ZN(n5237)
         );
  OAI22_X1 U2200 ( .A1(n3088), .A2(n3566), .B1(n3269), .B2(n2890), .ZN(n5238)
         );
  OAI22_X1 U2201 ( .A1(n3079), .A2(n3566), .B1(n3269), .B2(n2889), .ZN(n5239)
         );
  OAI22_X1 U2202 ( .A1(n3141), .A2(n3567), .B1(n7217), .B2(n2888), .ZN(n5240)
         );
  OAI22_X1 U2203 ( .A1(n3133), .A2(n3567), .B1(n7217), .B2(n2887), .ZN(n5241)
         );
  OAI22_X1 U2204 ( .A1(n3123), .A2(n3567), .B1(n7217), .B2(n2886), .ZN(n5242)
         );
  OAI22_X1 U2205 ( .A1(n3115), .A2(n3567), .B1(n7217), .B2(n2885), .ZN(n5243)
         );
  OAI22_X1 U2206 ( .A1(n3104), .A2(n3567), .B1(n7217), .B2(n2884), .ZN(n5244)
         );
  OAI22_X1 U2207 ( .A1(n3097), .A2(n3567), .B1(n7217), .B2(n2883), .ZN(n5245)
         );
  OAI22_X1 U2208 ( .A1(n3089), .A2(n3567), .B1(n7217), .B2(n2882), .ZN(n5246)
         );
  OAI22_X1 U2209 ( .A1(n3080), .A2(n3567), .B1(n7217), .B2(n2881), .ZN(n5247)
         );
  OAI22_X1 U2210 ( .A1(n3141), .A2(n3568), .B1(n3333), .B2(n2880), .ZN(n5248)
         );
  OAI22_X1 U2211 ( .A1(n3132), .A2(n3568), .B1(n3333), .B2(n2879), .ZN(n5249)
         );
  OAI22_X1 U2212 ( .A1(n3123), .A2(n3568), .B1(n3333), .B2(n2878), .ZN(n5250)
         );
  OAI22_X1 U2213 ( .A1(n3115), .A2(n3568), .B1(n3333), .B2(n2877), .ZN(n5251)
         );
  OAI22_X1 U2214 ( .A1(n3104), .A2(n3568), .B1(n3333), .B2(n2876), .ZN(n5252)
         );
  OAI22_X1 U2215 ( .A1(n3097), .A2(n3568), .B1(n3333), .B2(n2875), .ZN(n5253)
         );
  OAI22_X1 U2216 ( .A1(n3089), .A2(n3568), .B1(n3333), .B2(n2874), .ZN(n5254)
         );
  OAI22_X1 U2217 ( .A1(n3080), .A2(n3568), .B1(n3333), .B2(n2873), .ZN(n5255)
         );
  OAI22_X1 U2218 ( .A1(n3141), .A2(n3569), .B1(n7153), .B2(n2872), .ZN(n5256)
         );
  OAI22_X1 U2219 ( .A1(n3131), .A2(n3569), .B1(n7153), .B2(n2871), .ZN(n5257)
         );
  OAI22_X1 U2220 ( .A1(n3123), .A2(n3569), .B1(n7153), .B2(n2870), .ZN(n5258)
         );
  OAI22_X1 U2221 ( .A1(n3115), .A2(n3569), .B1(n7153), .B2(n2869), .ZN(n5259)
         );
  OAI22_X1 U2222 ( .A1(n3104), .A2(n3569), .B1(n7153), .B2(n2868), .ZN(n5260)
         );
  OAI22_X1 U2223 ( .A1(n3097), .A2(n3569), .B1(n7153), .B2(n2867), .ZN(n5261)
         );
  OAI22_X1 U2224 ( .A1(n3089), .A2(n3569), .B1(n7153), .B2(n2866), .ZN(n5262)
         );
  OAI22_X1 U2225 ( .A1(n3080), .A2(n3569), .B1(n7153), .B2(n2865), .ZN(n5263)
         );
  OAI22_X1 U2226 ( .A1(n3141), .A2(n3570), .B1(n3253), .B2(n2864), .ZN(n5264)
         );
  OAI22_X1 U2227 ( .A1(n3135), .A2(n3570), .B1(n3253), .B2(n2863), .ZN(n5265)
         );
  OAI22_X1 U2228 ( .A1(n3123), .A2(n3570), .B1(n3253), .B2(n2862), .ZN(n5266)
         );
  OAI22_X1 U2229 ( .A1(n3115), .A2(n3570), .B1(n3253), .B2(n2861), .ZN(n5267)
         );
  OAI22_X1 U2230 ( .A1(n3104), .A2(n3570), .B1(n3253), .B2(n2860), .ZN(n5268)
         );
  OAI22_X1 U2231 ( .A1(n3097), .A2(n3570), .B1(n3253), .B2(n2859), .ZN(n5269)
         );
  OAI22_X1 U2232 ( .A1(n3089), .A2(n3570), .B1(n3253), .B2(n2858), .ZN(n5270)
         );
  OAI22_X1 U2233 ( .A1(n3080), .A2(n3570), .B1(n3253), .B2(n2857), .ZN(n5271)
         );
  OAI22_X1 U2234 ( .A1(n3141), .A2(n3571), .B1(n7201), .B2(n2856), .ZN(n5272)
         );
  OAI22_X1 U2235 ( .A1(n3136), .A2(n3571), .B1(n7201), .B2(n2855), .ZN(n5273)
         );
  OAI22_X1 U2236 ( .A1(n3123), .A2(n3571), .B1(n7201), .B2(n2854), .ZN(n5274)
         );
  OAI22_X1 U2237 ( .A1(n3115), .A2(n3571), .B1(n7201), .B2(n2853), .ZN(n5275)
         );
  OAI22_X1 U2238 ( .A1(n3104), .A2(n3571), .B1(n7201), .B2(n2852), .ZN(n5276)
         );
  OAI22_X1 U2239 ( .A1(n3097), .A2(n3571), .B1(n7201), .B2(n2851), .ZN(n5277)
         );
  OAI22_X1 U2240 ( .A1(n3089), .A2(n3571), .B1(n7201), .B2(n2850), .ZN(n5278)
         );
  OAI22_X1 U2241 ( .A1(n3080), .A2(n3571), .B1(n7201), .B2(n2849), .ZN(n5279)
         );
  OAI22_X1 U2242 ( .A1(n3141), .A2(n3572), .B1(n3317), .B2(n2848), .ZN(n5280)
         );
  OAI22_X1 U2243 ( .A1(n3135), .A2(n3572), .B1(n3317), .B2(n2847), .ZN(n5281)
         );
  OAI22_X1 U2244 ( .A1(n3123), .A2(n3572), .B1(n3317), .B2(n2846), .ZN(n5282)
         );
  OAI22_X1 U2245 ( .A1(n3115), .A2(n3572), .B1(n3317), .B2(n2845), .ZN(n5283)
         );
  OAI22_X1 U2246 ( .A1(n3104), .A2(n3572), .B1(n3317), .B2(n2844), .ZN(n5284)
         );
  OAI22_X1 U2247 ( .A1(n3097), .A2(n3572), .B1(n3317), .B2(n2843), .ZN(n5285)
         );
  OAI22_X1 U2248 ( .A1(n3089), .A2(n3572), .B1(n3317), .B2(n2842), .ZN(n5286)
         );
  OAI22_X1 U2249 ( .A1(n3080), .A2(n3572), .B1(n3317), .B2(n2841), .ZN(n5287)
         );
  OAI22_X1 U2250 ( .A1(n3141), .A2(n3573), .B1(n7137), .B2(n2840), .ZN(n5288)
         );
  OAI22_X1 U2251 ( .A1(n3136), .A2(n3573), .B1(n7137), .B2(n2839), .ZN(n5289)
         );
  OAI22_X1 U2252 ( .A1(n3123), .A2(n3573), .B1(n7137), .B2(n2838), .ZN(n5290)
         );
  OAI22_X1 U2253 ( .A1(n3115), .A2(n3573), .B1(n7137), .B2(n2837), .ZN(n5291)
         );
  OAI22_X1 U2254 ( .A1(n3104), .A2(n3573), .B1(n7137), .B2(n2836), .ZN(n5292)
         );
  OAI22_X1 U2255 ( .A1(n3097), .A2(n3573), .B1(n7137), .B2(n2835), .ZN(n5293)
         );
  OAI22_X1 U2256 ( .A1(n3089), .A2(n3573), .B1(n7137), .B2(n2834), .ZN(n5294)
         );
  OAI22_X1 U2257 ( .A1(n3080), .A2(n3573), .B1(n7137), .B2(n2833), .ZN(n5295)
         );
  OAI22_X1 U2258 ( .A1(n3140), .A2(n3574), .B1(n3237), .B2(n2832), .ZN(n5296)
         );
  OAI22_X1 U2259 ( .A1(n3131), .A2(n3574), .B1(n3237), .B2(n2831), .ZN(n5297)
         );
  OAI22_X1 U2260 ( .A1(n3123), .A2(n3574), .B1(n3237), .B2(n2830), .ZN(n5298)
         );
  OAI22_X1 U2261 ( .A1(n3115), .A2(n3574), .B1(n3237), .B2(n2829), .ZN(n5299)
         );
  OAI22_X1 U2262 ( .A1(n3104), .A2(n3574), .B1(n3237), .B2(n2828), .ZN(n5300)
         );
  OAI22_X1 U2263 ( .A1(n3097), .A2(n3574), .B1(n3237), .B2(n2827), .ZN(n5301)
         );
  OAI22_X1 U2264 ( .A1(n3089), .A2(n3574), .B1(n3237), .B2(n2826), .ZN(n5302)
         );
  OAI22_X1 U2265 ( .A1(n3080), .A2(n3574), .B1(n3237), .B2(n2825), .ZN(n5303)
         );
  OAI22_X1 U2266 ( .A1(n3140), .A2(n3575), .B1(n7185), .B2(n2824), .ZN(n5304)
         );
  OAI22_X1 U2267 ( .A1(n3134), .A2(n3575), .B1(n7185), .B2(n2823), .ZN(n5305)
         );
  OAI22_X1 U2268 ( .A1(n3124), .A2(n3575), .B1(n7185), .B2(n2822), .ZN(n5306)
         );
  OAI22_X1 U2269 ( .A1(n3115), .A2(n3575), .B1(n7185), .B2(n2821), .ZN(n5307)
         );
  OAI22_X1 U2270 ( .A1(n3104), .A2(n3575), .B1(n7185), .B2(n2820), .ZN(n5308)
         );
  OAI22_X1 U2271 ( .A1(n3097), .A2(n3575), .B1(n7185), .B2(n2819), .ZN(n5309)
         );
  OAI22_X1 U2272 ( .A1(n3089), .A2(n3575), .B1(n7185), .B2(n2818), .ZN(n5310)
         );
  OAI22_X1 U2273 ( .A1(n3080), .A2(n3575), .B1(n7185), .B2(n2817), .ZN(n5311)
         );
  OAI22_X1 U2274 ( .A1(n3140), .A2(n3576), .B1(n3301), .B2(n2816), .ZN(n5312)
         );
  OAI22_X1 U2275 ( .A1(n3133), .A2(n3576), .B1(n3301), .B2(n2815), .ZN(n5313)
         );
  OAI22_X1 U2276 ( .A1(n3123), .A2(n3576), .B1(n3301), .B2(n2814), .ZN(n5314)
         );
  OAI22_X1 U2277 ( .A1(n3115), .A2(n3576), .B1(n3301), .B2(n2813), .ZN(n5315)
         );
  OAI22_X1 U2278 ( .A1(n3104), .A2(n3576), .B1(n3301), .B2(n2812), .ZN(n5316)
         );
  OAI22_X1 U2279 ( .A1(n3097), .A2(n3576), .B1(n3301), .B2(n2811), .ZN(n5317)
         );
  OAI22_X1 U2280 ( .A1(n3089), .A2(n3576), .B1(n3301), .B2(n2810), .ZN(n5318)
         );
  OAI22_X1 U2281 ( .A1(n3080), .A2(n3576), .B1(n3301), .B2(n2809), .ZN(n5319)
         );
  OAI22_X1 U2282 ( .A1(n3140), .A2(n3578), .B1(n7121), .B2(n2808), .ZN(n5320)
         );
  OAI22_X1 U2283 ( .A1(n3132), .A2(n3578), .B1(n7121), .B2(n2807), .ZN(n5321)
         );
  OAI22_X1 U2284 ( .A1(n3124), .A2(n3578), .B1(n7121), .B2(n2806), .ZN(n5322)
         );
  OAI22_X1 U2285 ( .A1(n3115), .A2(n3578), .B1(n7121), .B2(n2805), .ZN(n5323)
         );
  OAI22_X1 U2286 ( .A1(n3104), .A2(n3578), .B1(n7121), .B2(n2804), .ZN(n5324)
         );
  OAI22_X1 U2287 ( .A1(n3097), .A2(n3578), .B1(n7121), .B2(n2803), .ZN(n5325)
         );
  OAI22_X1 U2288 ( .A1(n3089), .A2(n3578), .B1(n7121), .B2(n2802), .ZN(n5326)
         );
  OAI22_X1 U2289 ( .A1(n3080), .A2(n3578), .B1(n7121), .B2(n2801), .ZN(n5327)
         );
  OAI22_X1 U2290 ( .A1(n3140), .A2(n3579), .B1(n3284), .B2(n2800), .ZN(n5328)
         );
  OAI22_X1 U2291 ( .A1(n3135), .A2(n3579), .B1(n3284), .B2(n2799), .ZN(n5329)
         );
  OAI22_X1 U2292 ( .A1(n3123), .A2(n3579), .B1(n3284), .B2(n2798), .ZN(n5330)
         );
  OAI22_X1 U2293 ( .A1(n3115), .A2(n3579), .B1(n3284), .B2(n2797), .ZN(n5331)
         );
  OAI22_X1 U2294 ( .A1(n3104), .A2(n3579), .B1(n3284), .B2(n2796), .ZN(n5332)
         );
  OAI22_X1 U2295 ( .A1(n3097), .A2(n3579), .B1(n3284), .B2(n2795), .ZN(n5333)
         );
  OAI22_X1 U2296 ( .A1(n3089), .A2(n3579), .B1(n3284), .B2(n2794), .ZN(n5334)
         );
  OAI22_X1 U2297 ( .A1(n3080), .A2(n3579), .B1(n3284), .B2(n2793), .ZN(n5335)
         );
  OAI22_X1 U2298 ( .A1(n3140), .A2(n3580), .B1(n7232), .B2(n2792), .ZN(n5336)
         );
  OAI22_X1 U2299 ( .A1(n3136), .A2(n3580), .B1(n7232), .B2(n2791), .ZN(n5337)
         );
  OAI22_X1 U2300 ( .A1(n3124), .A2(n3580), .B1(n7232), .B2(n2790), .ZN(n5338)
         );
  OAI22_X1 U2301 ( .A1(n3115), .A2(n3580), .B1(n7232), .B2(n2789), .ZN(n5339)
         );
  OAI22_X1 U2302 ( .A1(n3104), .A2(n3580), .B1(n7232), .B2(n2788), .ZN(n5340)
         );
  OAI22_X1 U2303 ( .A1(n3097), .A2(n3580), .B1(n7232), .B2(n2787), .ZN(n5341)
         );
  OAI22_X1 U2304 ( .A1(n3089), .A2(n3580), .B1(n7232), .B2(n2786), .ZN(n5342)
         );
  OAI22_X1 U2305 ( .A1(n3080), .A2(n3580), .B1(n7232), .B2(n2785), .ZN(n5343)
         );
  OAI22_X1 U2306 ( .A1(n3140), .A2(n3581), .B1(n3348), .B2(n2784), .ZN(n5344)
         );
  OAI22_X1 U2307 ( .A1(n3131), .A2(n3581), .B1(n3348), .B2(n2783), .ZN(n5345)
         );
  OAI22_X1 U2308 ( .A1(n3123), .A2(n3581), .B1(n3348), .B2(n2782), .ZN(n5346)
         );
  OAI22_X1 U2309 ( .A1(n3112), .A2(n3581), .B1(n3348), .B2(n2781), .ZN(n5347)
         );
  OAI22_X1 U2310 ( .A1(n3105), .A2(n3581), .B1(n3348), .B2(n2780), .ZN(n5348)
         );
  OAI22_X1 U2311 ( .A1(n3098), .A2(n3581), .B1(n3348), .B2(n2779), .ZN(n5349)
         );
  OAI22_X1 U2312 ( .A1(n3082), .A2(n3581), .B1(n3348), .B2(n2778), .ZN(n5350)
         );
  OAI22_X1 U2313 ( .A1(n3073), .A2(n3581), .B1(n3348), .B2(n2777), .ZN(n5351)
         );
  OAI22_X1 U2314 ( .A1(n3140), .A2(n3582), .B1(n7168), .B2(n2776), .ZN(n5352)
         );
  OAI22_X1 U2315 ( .A1(n3133), .A2(n3582), .B1(n7168), .B2(n2775), .ZN(n5353)
         );
  OAI22_X1 U2316 ( .A1(n3124), .A2(n3582), .B1(n7168), .B2(n2774), .ZN(n5354)
         );
  OAI22_X1 U2317 ( .A1(n3109), .A2(n3582), .B1(n7168), .B2(n2773), .ZN(n5355)
         );
  OAI22_X1 U2318 ( .A1(n3105), .A2(n3582), .B1(n7168), .B2(n2772), .ZN(n5356)
         );
  OAI22_X1 U2319 ( .A1(n3098), .A2(n3582), .B1(n7168), .B2(n2771), .ZN(n5357)
         );
  OAI22_X1 U2320 ( .A1(n3082), .A2(n3582), .B1(n7168), .B2(n2770), .ZN(n5358)
         );
  OAI22_X1 U2321 ( .A1(n3073), .A2(n3582), .B1(n7168), .B2(n2769), .ZN(n5359)
         );
  OAI22_X1 U2322 ( .A1(n3140), .A2(n3583), .B1(n3268), .B2(n2768), .ZN(n5360)
         );
  OAI22_X1 U2323 ( .A1(n3134), .A2(n3583), .B1(n3268), .B2(n2767), .ZN(n5361)
         );
  OAI22_X1 U2324 ( .A1(n3123), .A2(n3583), .B1(n3268), .B2(n2766), .ZN(n5362)
         );
  OAI22_X1 U2325 ( .A1(n3113), .A2(n3583), .B1(n3268), .B2(n2765), .ZN(n5363)
         );
  OAI22_X1 U2326 ( .A1(n3105), .A2(n3583), .B1(n3268), .B2(n2764), .ZN(n5364)
         );
  OAI22_X1 U2327 ( .A1(n3098), .A2(n3583), .B1(n3268), .B2(n2763), .ZN(n5365)
         );
  OAI22_X1 U2328 ( .A1(n3083), .A2(n3583), .B1(n3268), .B2(n2762), .ZN(n5366)
         );
  OAI22_X1 U2329 ( .A1(n3074), .A2(n3583), .B1(n3268), .B2(n2761), .ZN(n5367)
         );
  OAI22_X1 U2330 ( .A1(n3140), .A2(n3584), .B1(n7216), .B2(n2760), .ZN(n5368)
         );
  OAI22_X1 U2331 ( .A1(n3132), .A2(n3584), .B1(n7216), .B2(n2759), .ZN(n5369)
         );
  OAI22_X1 U2332 ( .A1(n3124), .A2(n3584), .B1(n7216), .B2(n2758), .ZN(n5370)
         );
  OAI22_X1 U2333 ( .A1(n3109), .A2(n3584), .B1(n7216), .B2(n2757), .ZN(n5371)
         );
  OAI22_X1 U2334 ( .A1(n3105), .A2(n3584), .B1(n7216), .B2(n2756), .ZN(n5372)
         );
  OAI22_X1 U2335 ( .A1(n3098), .A2(n3584), .B1(n7216), .B2(n2755), .ZN(n5373)
         );
  OAI22_X1 U2336 ( .A1(n3083), .A2(n3584), .B1(n7216), .B2(n2754), .ZN(n5374)
         );
  OAI22_X1 U2337 ( .A1(n3074), .A2(n3584), .B1(n7216), .B2(n2753), .ZN(n5375)
         );
  OAI22_X1 U2338 ( .A1(n3140), .A2(n3585), .B1(n3332), .B2(n2752), .ZN(n5376)
         );
  OAI22_X1 U2339 ( .A1(n3135), .A2(n3585), .B1(n3332), .B2(n2751), .ZN(n5377)
         );
  OAI22_X1 U2340 ( .A1(n3123), .A2(n3585), .B1(n3332), .B2(n2750), .ZN(n5378)
         );
  OAI22_X1 U2341 ( .A1(n3113), .A2(n3585), .B1(n3332), .B2(n2749), .ZN(n5379)
         );
  OAI22_X1 U2342 ( .A1(n3105), .A2(n3585), .B1(n3332), .B2(n2748), .ZN(n5380)
         );
  OAI22_X1 U2343 ( .A1(n3098), .A2(n3585), .B1(n3332), .B2(n2747), .ZN(n5381)
         );
  OAI22_X1 U2344 ( .A1(n3083), .A2(n3585), .B1(n3332), .B2(n2746), .ZN(n5382)
         );
  OAI22_X1 U2345 ( .A1(n3074), .A2(n3585), .B1(n3332), .B2(n2745), .ZN(n5383)
         );
  OAI22_X1 U2346 ( .A1(n3140), .A2(n3586), .B1(n7152), .B2(n2744), .ZN(n5384)
         );
  OAI22_X1 U2347 ( .A1(n3136), .A2(n3586), .B1(n7152), .B2(n2743), .ZN(n5385)
         );
  OAI22_X1 U2348 ( .A1(n3124), .A2(n3586), .B1(n7152), .B2(n2742), .ZN(n5386)
         );
  OAI22_X1 U2349 ( .A1(n3109), .A2(n3586), .B1(n7152), .B2(n2741), .ZN(n5387)
         );
  OAI22_X1 U2350 ( .A1(n3105), .A2(n3586), .B1(n7152), .B2(n2740), .ZN(n5388)
         );
  OAI22_X1 U2351 ( .A1(n3098), .A2(n3586), .B1(n7152), .B2(n2739), .ZN(n5389)
         );
  OAI22_X1 U2352 ( .A1(n3082), .A2(n3586), .B1(n7152), .B2(n2738), .ZN(n5390)
         );
  OAI22_X1 U2353 ( .A1(n3073), .A2(n3586), .B1(n7152), .B2(n2737), .ZN(n5391)
         );
  OAI22_X1 U2354 ( .A1(n3138), .A2(n3587), .B1(n3252), .B2(n2736), .ZN(n5392)
         );
  OAI22_X1 U2355 ( .A1(n3134), .A2(n3587), .B1(n3252), .B2(n2735), .ZN(n5393)
         );
  OAI22_X1 U2356 ( .A1(n3122), .A2(n3587), .B1(n3252), .B2(n2734), .ZN(n5394)
         );
  OAI22_X1 U2357 ( .A1(n3114), .A2(n3587), .B1(n3252), .B2(n2733), .ZN(n5395)
         );
  OAI22_X1 U2358 ( .A1(n3105), .A2(n3587), .B1(n3252), .B2(n2732), .ZN(n5396)
         );
  OAI22_X1 U2359 ( .A1(n3098), .A2(n3587), .B1(n3252), .B2(n2731), .ZN(n5397)
         );
  OAI22_X1 U2360 ( .A1(n3082), .A2(n3587), .B1(n3252), .B2(n2730), .ZN(n5398)
         );
  OAI22_X1 U2361 ( .A1(n3073), .A2(n3587), .B1(n3252), .B2(n2729), .ZN(n5399)
         );
  OAI22_X1 U2362 ( .A1(n3138), .A2(n3588), .B1(n7200), .B2(n2728), .ZN(n5400)
         );
  OAI22_X1 U2363 ( .A1(n3134), .A2(n3588), .B1(n7200), .B2(n2727), .ZN(n5401)
         );
  OAI22_X1 U2364 ( .A1(n3122), .A2(n3588), .B1(n7200), .B2(n2726), .ZN(n5402)
         );
  OAI22_X1 U2365 ( .A1(n3109), .A2(n3588), .B1(n7200), .B2(n2725), .ZN(n5403)
         );
  OAI22_X1 U2366 ( .A1(n3105), .A2(n3588), .B1(n7200), .B2(n2724), .ZN(n5404)
         );
  OAI22_X1 U2367 ( .A1(n3098), .A2(n3588), .B1(n7200), .B2(n2723), .ZN(n5405)
         );
  OAI22_X1 U2368 ( .A1(n3082), .A2(n3588), .B1(n7200), .B2(n2722), .ZN(n5406)
         );
  OAI22_X1 U2369 ( .A1(n3073), .A2(n3588), .B1(n7200), .B2(n2721), .ZN(n5407)
         );
  OAI22_X1 U2370 ( .A1(n3142), .A2(n3589), .B1(n3316), .B2(n2720), .ZN(n5408)
         );
  OAI22_X1 U2371 ( .A1(n3134), .A2(n3589), .B1(n3316), .B2(n2719), .ZN(n5409)
         );
  OAI22_X1 U2372 ( .A1(n3122), .A2(n3589), .B1(n3316), .B2(n2718), .ZN(n5410)
         );
  OAI22_X1 U2373 ( .A1(n3115), .A2(n3589), .B1(n3316), .B2(n2717), .ZN(n5411)
         );
  OAI22_X1 U2374 ( .A1(n3105), .A2(n3589), .B1(n3316), .B2(n2716), .ZN(n5412)
         );
  OAI22_X1 U2375 ( .A1(n3098), .A2(n3589), .B1(n3316), .B2(n2715), .ZN(n5413)
         );
  OAI22_X1 U2376 ( .A1(n3082), .A2(n3589), .B1(n3316), .B2(n2714), .ZN(n5414)
         );
  OAI22_X1 U2377 ( .A1(n3073), .A2(n3589), .B1(n3316), .B2(n2713), .ZN(n5415)
         );
  OAI22_X1 U2378 ( .A1(n3141), .A2(n3590), .B1(n7136), .B2(n2712), .ZN(n5416)
         );
  OAI22_X1 U2379 ( .A1(n3134), .A2(n3590), .B1(n7136), .B2(n2711), .ZN(n5417)
         );
  OAI22_X1 U2380 ( .A1(n3122), .A2(n3590), .B1(n7136), .B2(n2710), .ZN(n5418)
         );
  OAI22_X1 U2381 ( .A1(n3109), .A2(n3590), .B1(n7136), .B2(n2709), .ZN(n5419)
         );
  OAI22_X1 U2382 ( .A1(n3105), .A2(n3590), .B1(n7136), .B2(n2708), .ZN(n5420)
         );
  OAI22_X1 U2383 ( .A1(n3098), .A2(n3590), .B1(n7136), .B2(n2707), .ZN(n5421)
         );
  OAI22_X1 U2384 ( .A1(n3082), .A2(n3590), .B1(n7136), .B2(n2706), .ZN(n5422)
         );
  OAI22_X1 U2385 ( .A1(n3073), .A2(n3590), .B1(n7136), .B2(n2705), .ZN(n5423)
         );
  OAI22_X1 U2386 ( .A1(n3145), .A2(n3591), .B1(n3236), .B2(n2704), .ZN(n5424)
         );
  OAI22_X1 U2387 ( .A1(n3134), .A2(n3591), .B1(n3236), .B2(n2703), .ZN(n5425)
         );
  OAI22_X1 U2388 ( .A1(n3122), .A2(n3591), .B1(n3236), .B2(n2702), .ZN(n5426)
         );
  OAI22_X1 U2389 ( .A1(n3112), .A2(n3591), .B1(n3236), .B2(n2701), .ZN(n5427)
         );
  OAI22_X1 U2390 ( .A1(n3105), .A2(n3591), .B1(n3236), .B2(n2700), .ZN(n5428)
         );
  OAI22_X1 U2391 ( .A1(n3098), .A2(n3591), .B1(n3236), .B2(n2699), .ZN(n5429)
         );
  OAI22_X1 U2392 ( .A1(n3082), .A2(n3591), .B1(n3236), .B2(n2698), .ZN(n5430)
         );
  OAI22_X1 U2393 ( .A1(n3073), .A2(n3591), .B1(n3236), .B2(n2697), .ZN(n5431)
         );
  OAI22_X1 U2394 ( .A1(n3138), .A2(n3592), .B1(n7184), .B2(n2696), .ZN(n5432)
         );
  OAI22_X1 U2395 ( .A1(n3134), .A2(n3592), .B1(n7184), .B2(n2695), .ZN(n5433)
         );
  OAI22_X1 U2396 ( .A1(n3122), .A2(n3592), .B1(n7184), .B2(n2694), .ZN(n5434)
         );
  OAI22_X1 U2397 ( .A1(n3109), .A2(n3592), .B1(n7184), .B2(n2693), .ZN(n5435)
         );
  OAI22_X1 U2398 ( .A1(n3105), .A2(n3592), .B1(n7184), .B2(n2692), .ZN(n5436)
         );
  OAI22_X1 U2399 ( .A1(n3098), .A2(n3592), .B1(n7184), .B2(n2691), .ZN(n5437)
         );
  OAI22_X1 U2400 ( .A1(n3082), .A2(n3592), .B1(n7184), .B2(n2690), .ZN(n5438)
         );
  OAI22_X1 U2401 ( .A1(n3073), .A2(n3592), .B1(n7184), .B2(n2689), .ZN(n5439)
         );
  OAI22_X1 U2402 ( .A1(n3142), .A2(n3593), .B1(n3300), .B2(n2688), .ZN(n5440)
         );
  OAI22_X1 U2403 ( .A1(n3134), .A2(n3593), .B1(n3300), .B2(n2687), .ZN(n5441)
         );
  OAI22_X1 U2404 ( .A1(n3122), .A2(n3593), .B1(n3300), .B2(n2686), .ZN(n5442)
         );
  OAI22_X1 U2405 ( .A1(n3113), .A2(n3593), .B1(n3300), .B2(n2685), .ZN(n5443)
         );
  OAI22_X1 U2406 ( .A1(n3105), .A2(n3593), .B1(n3300), .B2(n2684), .ZN(n5444)
         );
  OAI22_X1 U2407 ( .A1(n3098), .A2(n3593), .B1(n3300), .B2(n2683), .ZN(n5445)
         );
  OAI22_X1 U2408 ( .A1(n3082), .A2(n3593), .B1(n3300), .B2(n2682), .ZN(n5446)
         );
  OAI22_X1 U2409 ( .A1(n3073), .A2(n3593), .B1(n3300), .B2(n2681), .ZN(n5447)
         );
  OAI22_X1 U2410 ( .A1(n3141), .A2(n3595), .B1(n7120), .B2(n2680), .ZN(n5448)
         );
  OAI22_X1 U2411 ( .A1(n3134), .A2(n3595), .B1(n7120), .B2(n2679), .ZN(n5449)
         );
  OAI22_X1 U2412 ( .A1(n3122), .A2(n3595), .B1(n7120), .B2(n2678), .ZN(n5450)
         );
  OAI22_X1 U2413 ( .A1(n3114), .A2(n3595), .B1(n7120), .B2(n2677), .ZN(n5451)
         );
  OAI22_X1 U2414 ( .A1(n3106), .A2(n3595), .B1(n7120), .B2(n2676), .ZN(n5452)
         );
  OAI22_X1 U2415 ( .A1(n3099), .A2(n3595), .B1(n7120), .B2(n2675), .ZN(n5453)
         );
  OAI22_X1 U2416 ( .A1(n3082), .A2(n3595), .B1(n7120), .B2(n2674), .ZN(n5454)
         );
  OAI22_X1 U2417 ( .A1(n3073), .A2(n3595), .B1(n7120), .B2(n2673), .ZN(n5455)
         );
  OAI22_X1 U2418 ( .A1(n3145), .A2(n3596), .B1(n3283), .B2(n2672), .ZN(n5456)
         );
  OAI22_X1 U2419 ( .A1(n3134), .A2(n3596), .B1(n3283), .B2(n2671), .ZN(n5457)
         );
  OAI22_X1 U2420 ( .A1(n3122), .A2(n3596), .B1(n3283), .B2(n2670), .ZN(n5458)
         );
  OAI22_X1 U2421 ( .A1(n3109), .A2(n3596), .B1(n3283), .B2(n2669), .ZN(n5459)
         );
  OAI22_X1 U2422 ( .A1(n3106), .A2(n3596), .B1(n3283), .B2(n2668), .ZN(n5460)
         );
  OAI22_X1 U2423 ( .A1(n3099), .A2(n3596), .B1(n3283), .B2(n2667), .ZN(n5461)
         );
  OAI22_X1 U2424 ( .A1(n3082), .A2(n3596), .B1(n3283), .B2(n2666), .ZN(n5462)
         );
  OAI22_X1 U2425 ( .A1(n3073), .A2(n3596), .B1(n3283), .B2(n2665), .ZN(n5463)
         );
  OAI22_X1 U2426 ( .A1(n3137), .A2(n3597), .B1(n7231), .B2(n2664), .ZN(n5464)
         );
  OAI22_X1 U2427 ( .A1(n3134), .A2(n3597), .B1(n7231), .B2(n2663), .ZN(n5465)
         );
  OAI22_X1 U2428 ( .A1(n3122), .A2(n3597), .B1(n7231), .B2(n2662), .ZN(n5466)
         );
  OAI22_X1 U2429 ( .A1(n3114), .A2(n3597), .B1(n7231), .B2(n2661), .ZN(n5467)
         );
  OAI22_X1 U2430 ( .A1(n3106), .A2(n3597), .B1(n7231), .B2(n2660), .ZN(n5468)
         );
  OAI22_X1 U2431 ( .A1(n3099), .A2(n3597), .B1(n7231), .B2(n2659), .ZN(n5469)
         );
  OAI22_X1 U2432 ( .A1(n3090), .A2(n3597), .B1(n7231), .B2(n2658), .ZN(n5470)
         );
  OAI22_X1 U2433 ( .A1(n3081), .A2(n3597), .B1(n7231), .B2(n2657), .ZN(n5471)
         );
  OAI22_X1 U2434 ( .A1(n3138), .A2(n3598), .B1(n3347), .B2(n2656), .ZN(n5472)
         );
  OAI22_X1 U2435 ( .A1(n3134), .A2(n3598), .B1(n3347), .B2(n2655), .ZN(n5473)
         );
  OAI22_X1 U2436 ( .A1(n3122), .A2(n3598), .B1(n3347), .B2(n2654), .ZN(n5474)
         );
  OAI22_X1 U2437 ( .A1(n3116), .A2(n3598), .B1(n3347), .B2(n2653), .ZN(n5475)
         );
  OAI22_X1 U2438 ( .A1(n3106), .A2(n3598), .B1(n3347), .B2(n2652), .ZN(n5476)
         );
  OAI22_X1 U2439 ( .A1(n3099), .A2(n3598), .B1(n3347), .B2(n2651), .ZN(n5477)
         );
  OAI22_X1 U2440 ( .A1(n3083), .A2(n3598), .B1(n3347), .B2(n2650), .ZN(n5478)
         );
  OAI22_X1 U2441 ( .A1(n3074), .A2(n3598), .B1(n3347), .B2(n2649), .ZN(n5479)
         );
  OAI22_X1 U2442 ( .A1(n3138), .A2(n3599), .B1(n7167), .B2(n2648), .ZN(n5480)
         );
  OAI22_X1 U2443 ( .A1(n3134), .A2(n3599), .B1(n7167), .B2(n2647), .ZN(n5481)
         );
  OAI22_X1 U2444 ( .A1(n3122), .A2(n3599), .B1(n7167), .B2(n2646), .ZN(n5482)
         );
  OAI22_X1 U2445 ( .A1(n3117), .A2(n3599), .B1(n7167), .B2(n2645), .ZN(n5483)
         );
  OAI22_X1 U2446 ( .A1(n3106), .A2(n3599), .B1(n7167), .B2(n2644), .ZN(n5484)
         );
  OAI22_X1 U2447 ( .A1(n3099), .A2(n3599), .B1(n7167), .B2(n2643), .ZN(n5485)
         );
  OAI22_X1 U2448 ( .A1(n3083), .A2(n3599), .B1(n7167), .B2(n2642), .ZN(n5486)
         );
  OAI22_X1 U2449 ( .A1(n3074), .A2(n3599), .B1(n7167), .B2(n2641), .ZN(n5487)
         );
  OAI22_X1 U2450 ( .A1(n3138), .A2(n3600), .B1(n3267), .B2(n2640), .ZN(n5488)
         );
  OAI22_X1 U2451 ( .A1(n3134), .A2(n3600), .B1(n3267), .B2(n2639), .ZN(n5489)
         );
  OAI22_X1 U2452 ( .A1(n3122), .A2(n3600), .B1(n3267), .B2(n2638), .ZN(n5490)
         );
  OAI22_X1 U2453 ( .A1(n3116), .A2(n3600), .B1(n3267), .B2(n2637), .ZN(n5491)
         );
  OAI22_X1 U2454 ( .A1(n3106), .A2(n3600), .B1(n3267), .B2(n2636), .ZN(n5492)
         );
  OAI22_X1 U2455 ( .A1(n3099), .A2(n3600), .B1(n3267), .B2(n2635), .ZN(n5493)
         );
  OAI22_X1 U2456 ( .A1(n3083), .A2(n3600), .B1(n3267), .B2(n2634), .ZN(n5494)
         );
  OAI22_X1 U2457 ( .A1(n3074), .A2(n3600), .B1(n3267), .B2(n2633), .ZN(n5495)
         );
  OAI22_X1 U2458 ( .A1(n3144), .A2(n3601), .B1(n7215), .B2(n2632), .ZN(n5496)
         );
  OAI22_X1 U2459 ( .A1(n3133), .A2(n3601), .B1(n7215), .B2(n2631), .ZN(n5497)
         );
  OAI22_X1 U2460 ( .A1(n3122), .A2(n3601), .B1(n7215), .B2(n2630), .ZN(n5498)
         );
  OAI22_X1 U2461 ( .A1(n3117), .A2(n3601), .B1(n7215), .B2(n2629), .ZN(n5499)
         );
  OAI22_X1 U2462 ( .A1(n3106), .A2(n3601), .B1(n7215), .B2(n2628), .ZN(n5500)
         );
  OAI22_X1 U2463 ( .A1(n3099), .A2(n3601), .B1(n7215), .B2(n2627), .ZN(n5501)
         );
  OAI22_X1 U2464 ( .A1(n3083), .A2(n3601), .B1(n7215), .B2(n2626), .ZN(n5502)
         );
  OAI22_X1 U2465 ( .A1(n3074), .A2(n3601), .B1(n7215), .B2(n2625), .ZN(n5503)
         );
  OAI22_X1 U2466 ( .A1(n3143), .A2(n3602), .B1(n3331), .B2(n2624), .ZN(n5504)
         );
  OAI22_X1 U2467 ( .A1(n3133), .A2(n3602), .B1(n3331), .B2(n2623), .ZN(n5505)
         );
  OAI22_X1 U2468 ( .A1(n3126), .A2(n3602), .B1(n3331), .B2(n2622), .ZN(n5506)
         );
  OAI22_X1 U2469 ( .A1(n3116), .A2(n3602), .B1(n3331), .B2(n2621), .ZN(n5507)
         );
  OAI22_X1 U2470 ( .A1(n3106), .A2(n3602), .B1(n3331), .B2(n2620), .ZN(n5508)
         );
  OAI22_X1 U2471 ( .A1(n3099), .A2(n3602), .B1(n3331), .B2(n2619), .ZN(n5509)
         );
  OAI22_X1 U2472 ( .A1(n3083), .A2(n3602), .B1(n3331), .B2(n2618), .ZN(n5510)
         );
  OAI22_X1 U2473 ( .A1(n3074), .A2(n3602), .B1(n3331), .B2(n2617), .ZN(n5511)
         );
  OAI22_X1 U2474 ( .A1(n3145), .A2(n3603), .B1(n7151), .B2(n2616), .ZN(n5512)
         );
  OAI22_X1 U2475 ( .A1(n3133), .A2(n3603), .B1(n7151), .B2(n2615), .ZN(n5513)
         );
  OAI22_X1 U2476 ( .A1(n3125), .A2(n3603), .B1(n7151), .B2(n2614), .ZN(n5514)
         );
  OAI22_X1 U2477 ( .A1(n3117), .A2(n3603), .B1(n7151), .B2(n2613), .ZN(n5515)
         );
  OAI22_X1 U2478 ( .A1(n3106), .A2(n3603), .B1(n7151), .B2(n2612), .ZN(n5516)
         );
  OAI22_X1 U2479 ( .A1(n3099), .A2(n3603), .B1(n7151), .B2(n2611), .ZN(n5517)
         );
  OAI22_X1 U2480 ( .A1(n3083), .A2(n3603), .B1(n7151), .B2(n2610), .ZN(n5518)
         );
  OAI22_X1 U2481 ( .A1(n3074), .A2(n3603), .B1(n7151), .B2(n2609), .ZN(n5519)
         );
  OAI22_X1 U2482 ( .A1(n3145), .A2(n3604), .B1(n3251), .B2(n2592), .ZN(n5520)
         );
  OAI22_X1 U2483 ( .A1(n3133), .A2(n3604), .B1(n3251), .B2(n2591), .ZN(n5521)
         );
  OAI22_X1 U2484 ( .A1(n3127), .A2(n3604), .B1(n3251), .B2(n2590), .ZN(n5522)
         );
  OAI22_X1 U2485 ( .A1(n3109), .A2(n3604), .B1(n3251), .B2(n2589), .ZN(n5523)
         );
  OAI22_X1 U2486 ( .A1(n3106), .A2(n3604), .B1(n3251), .B2(n2588), .ZN(n5524)
         );
  OAI22_X1 U2487 ( .A1(n3099), .A2(n3604), .B1(n3251), .B2(n2587), .ZN(n5525)
         );
  OAI22_X1 U2488 ( .A1(n3083), .A2(n3604), .B1(n3251), .B2(n2586), .ZN(n5526)
         );
  OAI22_X1 U2489 ( .A1(n3074), .A2(n3604), .B1(n3251), .B2(n2585), .ZN(n5527)
         );
  OAI22_X1 U2490 ( .A1(n3138), .A2(n3605), .B1(n7199), .B2(n2584), .ZN(n5528)
         );
  OAI22_X1 U2491 ( .A1(n3133), .A2(n3605), .B1(n7199), .B2(n2583), .ZN(n5529)
         );
  OAI22_X1 U2492 ( .A1(n3122), .A2(n3605), .B1(n7199), .B2(n2582), .ZN(n5530)
         );
  OAI22_X1 U2493 ( .A1(n3115), .A2(n3605), .B1(n7199), .B2(n2581), .ZN(n5531)
         );
  OAI22_X1 U2494 ( .A1(n3106), .A2(n3605), .B1(n7199), .B2(n2580), .ZN(n5532)
         );
  OAI22_X1 U2495 ( .A1(n3099), .A2(n3605), .B1(n7199), .B2(n2579), .ZN(n5533)
         );
  OAI22_X1 U2496 ( .A1(n3083), .A2(n3605), .B1(n7199), .B2(n2578), .ZN(n5534)
         );
  OAI22_X1 U2497 ( .A1(n3074), .A2(n3605), .B1(n7199), .B2(n2577), .ZN(n5535)
         );
  OAI22_X1 U2498 ( .A1(n3138), .A2(n3606), .B1(n3315), .B2(n2560), .ZN(n5536)
         );
  OAI22_X1 U2499 ( .A1(n3133), .A2(n3606), .B1(n3315), .B2(n2559), .ZN(n5537)
         );
  OAI22_X1 U2500 ( .A1(n3126), .A2(n3606), .B1(n3315), .B2(n2558), .ZN(n5538)
         );
  OAI22_X1 U2501 ( .A1(n3109), .A2(n3606), .B1(n3315), .B2(n2557), .ZN(n5539)
         );
  OAI22_X1 U2502 ( .A1(n3106), .A2(n3606), .B1(n3315), .B2(n2556), .ZN(n5540)
         );
  OAI22_X1 U2503 ( .A1(n3099), .A2(n3606), .B1(n3315), .B2(n2555), .ZN(n5541)
         );
  OAI22_X1 U2504 ( .A1(n3083), .A2(n3606), .B1(n3315), .B2(n2554), .ZN(n5542)
         );
  OAI22_X1 U2505 ( .A1(n3074), .A2(n3606), .B1(n3315), .B2(n2553), .ZN(n5543)
         );
  OAI22_X1 U2506 ( .A1(n3141), .A2(n3607), .B1(n7135), .B2(n2552), .ZN(n5544)
         );
  OAI22_X1 U2507 ( .A1(n3133), .A2(n3607), .B1(n7135), .B2(n2551), .ZN(n5545)
         );
  OAI22_X1 U2508 ( .A1(n3125), .A2(n3607), .B1(n7135), .B2(n2550), .ZN(n5546)
         );
  OAI22_X1 U2509 ( .A1(n3112), .A2(n3607), .B1(n7135), .B2(n2549), .ZN(n5547)
         );
  OAI22_X1 U2510 ( .A1(n3106), .A2(n3607), .B1(n7135), .B2(n2548), .ZN(n5548)
         );
  OAI22_X1 U2511 ( .A1(n3099), .A2(n3607), .B1(n7135), .B2(n2547), .ZN(n5549)
         );
  OAI22_X1 U2512 ( .A1(n3083), .A2(n3607), .B1(n7135), .B2(n2546), .ZN(n5550)
         );
  OAI22_X1 U2513 ( .A1(n3074), .A2(n3607), .B1(n7135), .B2(n2545), .ZN(n5551)
         );
  OAI22_X1 U2514 ( .A1(n3144), .A2(n3608), .B1(n3235), .B2(n2528), .ZN(n5552)
         );
  OAI22_X1 U2515 ( .A1(n3133), .A2(n3608), .B1(n3235), .B2(n2527), .ZN(n5553)
         );
  OAI22_X1 U2516 ( .A1(n3127), .A2(n3608), .B1(n3235), .B2(n2526), .ZN(n5554)
         );
  OAI22_X1 U2517 ( .A1(n3113), .A2(n3608), .B1(n3235), .B2(n2525), .ZN(n5555)
         );
  OAI22_X1 U2518 ( .A1(n3107), .A2(n3608), .B1(n3235), .B2(n2524), .ZN(n5556)
         );
  OAI22_X1 U2519 ( .A1(n3099), .A2(n3608), .B1(n3235), .B2(n2523), .ZN(n5557)
         );
  OAI22_X1 U2520 ( .A1(n3082), .A2(n3608), .B1(n3235), .B2(n2522), .ZN(n5558)
         );
  OAI22_X1 U2521 ( .A1(n3073), .A2(n3608), .B1(n3235), .B2(n2521), .ZN(n5559)
         );
  OAI22_X1 U2522 ( .A1(n3143), .A2(n3609), .B1(n7183), .B2(n2520), .ZN(n5560)
         );
  OAI22_X1 U2523 ( .A1(n3133), .A2(n3609), .B1(n7183), .B2(n2519), .ZN(n5561)
         );
  OAI22_X1 U2524 ( .A1(n3122), .A2(n3609), .B1(n7183), .B2(n2518), .ZN(n5562)
         );
  OAI22_X1 U2525 ( .A1(n3115), .A2(n3609), .B1(n7183), .B2(n2517), .ZN(n5563)
         );
  OAI22_X1 U2526 ( .A1(n3107), .A2(n3609), .B1(n7183), .B2(n2516), .ZN(n5564)
         );
  OAI22_X1 U2527 ( .A1(n3098), .A2(n3609), .B1(n7183), .B2(n2515), .ZN(n5565)
         );
  OAI22_X1 U2528 ( .A1(n3082), .A2(n3609), .B1(n7183), .B2(n2514), .ZN(n5566)
         );
  OAI22_X1 U2529 ( .A1(n3073), .A2(n3609), .B1(n7183), .B2(n2513), .ZN(n5567)
         );
  OAI22_X1 U2530 ( .A1(n3138), .A2(n3610), .B1(n3299), .B2(n2496), .ZN(n5568)
         );
  OAI22_X1 U2531 ( .A1(n3133), .A2(n3610), .B1(n3299), .B2(n2495), .ZN(n5569)
         );
  OAI22_X1 U2532 ( .A1(n3126), .A2(n3610), .B1(n3299), .B2(n2494), .ZN(n5570)
         );
  OAI22_X1 U2533 ( .A1(n3109), .A2(n3610), .B1(n3299), .B2(n2493), .ZN(n5571)
         );
  OAI22_X1 U2534 ( .A1(n3107), .A2(n3610), .B1(n3299), .B2(n2492), .ZN(n5572)
         );
  OAI22_X1 U2535 ( .A1(n3095), .A2(n3610), .B1(n3299), .B2(n2491), .ZN(n5573)
         );
  OAI22_X1 U2536 ( .A1(n3082), .A2(n3610), .B1(n3299), .B2(n2490), .ZN(n5574)
         );
  OAI22_X1 U2537 ( .A1(n3073), .A2(n3610), .B1(n3299), .B2(n2489), .ZN(n5575)
         );
  OAI22_X1 U2538 ( .A1(n3137), .A2(n3612), .B1(n7119), .B2(n2488), .ZN(n5576)
         );
  OAI22_X1 U2539 ( .A1(n3133), .A2(n3612), .B1(n7119), .B2(n2487), .ZN(n5577)
         );
  OAI22_X1 U2540 ( .A1(n3125), .A2(n3612), .B1(n7119), .B2(n2486), .ZN(n5578)
         );
  OAI22_X1 U2541 ( .A1(n3116), .A2(n3612), .B1(n7119), .B2(n2485), .ZN(n5579)
         );
  OAI22_X1 U2542 ( .A1(n3107), .A2(n3612), .B1(n7119), .B2(n2484), .ZN(n5580)
         );
  OAI22_X1 U2543 ( .A1(n3096), .A2(n3612), .B1(n7119), .B2(n2483), .ZN(n5581)
         );
  OAI22_X1 U2544 ( .A1(n3082), .A2(n3612), .B1(n7119), .B2(n2482), .ZN(n5582)
         );
  OAI22_X1 U2545 ( .A1(n3073), .A2(n3612), .B1(n7119), .B2(n2481), .ZN(n5583)
         );
  OAI22_X1 U2546 ( .A1(n3138), .A2(n3613), .B1(n3282), .B2(n2464), .ZN(n5584)
         );
  OAI22_X1 U2547 ( .A1(n3133), .A2(n3613), .B1(n3282), .B2(n2463), .ZN(n5585)
         );
  OAI22_X1 U2548 ( .A1(n3127), .A2(n3613), .B1(n3282), .B2(n2462), .ZN(n5586)
         );
  OAI22_X1 U2549 ( .A1(n3117), .A2(n3613), .B1(n3282), .B2(n2461), .ZN(n5587)
         );
  OAI22_X1 U2550 ( .A1(n3107), .A2(n3613), .B1(n3282), .B2(n2460), .ZN(n5588)
         );
  OAI22_X1 U2551 ( .A1(n3097), .A2(n3613), .B1(n3282), .B2(n2459), .ZN(n5589)
         );
  OAI22_X1 U2552 ( .A1(n3082), .A2(n3613), .B1(n3282), .B2(n2458), .ZN(n5590)
         );
  OAI22_X1 U2553 ( .A1(n3073), .A2(n3613), .B1(n3282), .B2(n2457), .ZN(n5591)
         );
  OAI22_X1 U2554 ( .A1(n3138), .A2(n3614), .B1(n7230), .B2(n2456), .ZN(n5592)
         );
  OAI22_X1 U2555 ( .A1(n3133), .A2(n3614), .B1(n7230), .B2(n2455), .ZN(n5593)
         );
  OAI22_X1 U2556 ( .A1(n3122), .A2(n3614), .B1(n7230), .B2(n2454), .ZN(n5594)
         );
  OAI22_X1 U2557 ( .A1(n3116), .A2(n3614), .B1(n7230), .B2(n2453), .ZN(n5595)
         );
  OAI22_X1 U2558 ( .A1(n3107), .A2(n3614), .B1(n7230), .B2(n2452), .ZN(n5596)
         );
  OAI22_X1 U2559 ( .A1(n3098), .A2(n3614), .B1(n7230), .B2(n2451), .ZN(n5597)
         );
  OAI22_X1 U2560 ( .A1(n3088), .A2(n3614), .B1(n7230), .B2(n2450), .ZN(n5598)
         );
  OAI22_X1 U2561 ( .A1(n3079), .A2(n3614), .B1(n7230), .B2(n2449), .ZN(n5599)
         );
  OAI22_X1 U2562 ( .A1(n3138), .A2(n3615), .B1(n3346), .B2(n2432), .ZN(n5600)
         );
  OAI22_X1 U2563 ( .A1(n3132), .A2(n3615), .B1(n3346), .B2(n2431), .ZN(n5601)
         );
  OAI22_X1 U2564 ( .A1(n3127), .A2(n3615), .B1(n3346), .B2(n2430), .ZN(n5602)
         );
  OAI22_X1 U2565 ( .A1(n3117), .A2(n3615), .B1(n3346), .B2(n2429), .ZN(n5603)
         );
  OAI22_X1 U2566 ( .A1(n3107), .A2(n3615), .B1(n3346), .B2(n2428), .ZN(n5604)
         );
  OAI22_X1 U2567 ( .A1(n3099), .A2(n3615), .B1(n3346), .B2(n2427), .ZN(n5605)
         );
  OAI22_X1 U2568 ( .A1(n3086), .A2(n3615), .B1(n3346), .B2(n2426), .ZN(n5606)
         );
  OAI22_X1 U2569 ( .A1(n3077), .A2(n3615), .B1(n3346), .B2(n2425), .ZN(n5607)
         );
  OAI22_X1 U2570 ( .A1(n3138), .A2(n3616), .B1(n7166), .B2(n2424), .ZN(n5608)
         );
  OAI22_X1 U2571 ( .A1(n3132), .A2(n3616), .B1(n7166), .B2(n2423), .ZN(n5609)
         );
  OAI22_X1 U2572 ( .A1(n3118), .A2(n3616), .B1(n7166), .B2(n2422), .ZN(n5610)
         );
  OAI22_X1 U2573 ( .A1(n3116), .A2(n3616), .B1(n7166), .B2(n2421), .ZN(n5611)
         );
  OAI22_X1 U2574 ( .A1(n3107), .A2(n3616), .B1(n7166), .B2(n2420), .ZN(n5612)
         );
  OAI22_X1 U2575 ( .A1(n3095), .A2(n3616), .B1(n7166), .B2(n2419), .ZN(n5613)
         );
  OAI22_X1 U2576 ( .A1(n3088), .A2(n3616), .B1(n7166), .B2(n2418), .ZN(n5614)
         );
  OAI22_X1 U2577 ( .A1(n3079), .A2(n3616), .B1(n7166), .B2(n2417), .ZN(n5615)
         );
  OAI22_X1 U2578 ( .A1(n3145), .A2(n3617), .B1(n3266), .B2(n2400), .ZN(n5616)
         );
  OAI22_X1 U2579 ( .A1(n3132), .A2(n3617), .B1(n3266), .B2(n2399), .ZN(n5617)
         );
  OAI22_X1 U2580 ( .A1(n3118), .A2(n3617), .B1(n3266), .B2(n2398), .ZN(n5618)
         );
  OAI22_X1 U2581 ( .A1(n3117), .A2(n3617), .B1(n3266), .B2(n2397), .ZN(n5619)
         );
  OAI22_X1 U2582 ( .A1(n3107), .A2(n3617), .B1(n3266), .B2(n2396), .ZN(n5620)
         );
  OAI22_X1 U2583 ( .A1(n3096), .A2(n3617), .B1(n3266), .B2(n2395), .ZN(n5621)
         );
  OAI22_X1 U2584 ( .A1(n3090), .A2(n3617), .B1(n3266), .B2(n2394), .ZN(n5622)
         );
  OAI22_X1 U2585 ( .A1(n3081), .A2(n3617), .B1(n3266), .B2(n2393), .ZN(n5623)
         );
  OAI22_X1 U2586 ( .A1(n3138), .A2(n3618), .B1(n7214), .B2(n2392), .ZN(n5624)
         );
  OAI22_X1 U2587 ( .A1(n3132), .A2(n3618), .B1(n7214), .B2(n2391), .ZN(n5625)
         );
  OAI22_X1 U2588 ( .A1(n3118), .A2(n3618), .B1(n7214), .B2(n2390), .ZN(n5626)
         );
  OAI22_X1 U2589 ( .A1(n3116), .A2(n3618), .B1(n7214), .B2(n2389), .ZN(n5627)
         );
  OAI22_X1 U2590 ( .A1(n3107), .A2(n3618), .B1(n7214), .B2(n2388), .ZN(n5628)
         );
  OAI22_X1 U2591 ( .A1(n3097), .A2(n3618), .B1(n7214), .B2(n2387), .ZN(n5629)
         );
  OAI22_X1 U2592 ( .A1(n3083), .A2(n3618), .B1(n7214), .B2(n2386), .ZN(n5630)
         );
  OAI22_X1 U2593 ( .A1(n3074), .A2(n3618), .B1(n7214), .B2(n2385), .ZN(n5631)
         );
  OAI22_X1 U2594 ( .A1(n3142), .A2(n3619), .B1(n3330), .B2(n2368), .ZN(n5632)
         );
  OAI22_X1 U2595 ( .A1(n3132), .A2(n3619), .B1(n3330), .B2(n2367), .ZN(n5633)
         );
  OAI22_X1 U2596 ( .A1(n3122), .A2(n3619), .B1(n3330), .B2(n2366), .ZN(n5634)
         );
  OAI22_X1 U2597 ( .A1(n3117), .A2(n3619), .B1(n3330), .B2(n2365), .ZN(n5635)
         );
  OAI22_X1 U2598 ( .A1(n3107), .A2(n3619), .B1(n3330), .B2(n2364), .ZN(n5636)
         );
  OAI22_X1 U2599 ( .A1(n3099), .A2(n3619), .B1(n3330), .B2(n2363), .ZN(n5637)
         );
  OAI22_X1 U2600 ( .A1(n3083), .A2(n3619), .B1(n3330), .B2(n2362), .ZN(n5638)
         );
  OAI22_X1 U2601 ( .A1(n3074), .A2(n3619), .B1(n3330), .B2(n2361), .ZN(n5639)
         );
  OAI22_X1 U2602 ( .A1(n3141), .A2(n3620), .B1(n7150), .B2(n2360), .ZN(n5640)
         );
  OAI22_X1 U2603 ( .A1(n3132), .A2(n3620), .B1(n7150), .B2(n2359), .ZN(n5641)
         );
  OAI22_X1 U2604 ( .A1(n3126), .A2(n3620), .B1(n7150), .B2(n2358), .ZN(n5642)
         );
  OAI22_X1 U2605 ( .A1(n3116), .A2(n3620), .B1(n7150), .B2(n2357), .ZN(n5643)
         );
  OAI22_X1 U2606 ( .A1(n3107), .A2(n3620), .B1(n7150), .B2(n2356), .ZN(n5644)
         );
  OAI22_X1 U2607 ( .A1(n3098), .A2(n3620), .B1(n7150), .B2(n2355), .ZN(n5645)
         );
  OAI22_X1 U2608 ( .A1(n3083), .A2(n3620), .B1(n7150), .B2(n2354), .ZN(n5646)
         );
  OAI22_X1 U2609 ( .A1(n3074), .A2(n3620), .B1(n7150), .B2(n2353), .ZN(n5647)
         );
  OAI22_X1 U2610 ( .A1(n3138), .A2(n3621), .B1(n3250), .B2(n2336), .ZN(n5648)
         );
  OAI22_X1 U2611 ( .A1(n3132), .A2(n3621), .B1(n3250), .B2(n2335), .ZN(n5649)
         );
  OAI22_X1 U2612 ( .A1(n3126), .A2(n3621), .B1(n3250), .B2(n2334), .ZN(n5650)
         );
  OAI22_X1 U2613 ( .A1(n3117), .A2(n3621), .B1(n3250), .B2(n2333), .ZN(n5651)
         );
  OAI22_X1 U2614 ( .A1(n3107), .A2(n3621), .B1(n3250), .B2(n2332), .ZN(n5652)
         );
  OAI22_X1 U2615 ( .A1(n3095), .A2(n3621), .B1(n3250), .B2(n2331), .ZN(n5653)
         );
  OAI22_X1 U2616 ( .A1(n3083), .A2(n3621), .B1(n3250), .B2(n2330), .ZN(n5654)
         );
  OAI22_X1 U2617 ( .A1(n3074), .A2(n3621), .B1(n3250), .B2(n2329), .ZN(n5655)
         );
  OAI22_X1 U2618 ( .A1(n3138), .A2(n3622), .B1(n7198), .B2(n2328), .ZN(n5656)
         );
  OAI22_X1 U2619 ( .A1(n3132), .A2(n3622), .B1(n7198), .B2(n2327), .ZN(n5657)
         );
  OAI22_X1 U2620 ( .A1(n3125), .A2(n3622), .B1(n7198), .B2(n2326), .ZN(n5658)
         );
  OAI22_X1 U2621 ( .A1(n3116), .A2(n3622), .B1(n7198), .B2(n2325), .ZN(n5659)
         );
  OAI22_X1 U2622 ( .A1(n3108), .A2(n3622), .B1(n7198), .B2(n2324), .ZN(n5660)
         );
  OAI22_X1 U2623 ( .A1(n3095), .A2(n3622), .B1(n7198), .B2(n2323), .ZN(n5661)
         );
  OAI22_X1 U2624 ( .A1(n3084), .A2(n3622), .B1(n7198), .B2(n2322), .ZN(n5662)
         );
  OAI22_X1 U2625 ( .A1(n3075), .A2(n3622), .B1(n7198), .B2(n2321), .ZN(n5663)
         );
  OAI22_X1 U2626 ( .A1(n3138), .A2(n3623), .B1(n3314), .B2(n2304), .ZN(n5664)
         );
  OAI22_X1 U2627 ( .A1(n3132), .A2(n3623), .B1(n3314), .B2(n2303), .ZN(n5665)
         );
  OAI22_X1 U2628 ( .A1(n3127), .A2(n3623), .B1(n3314), .B2(n2302), .ZN(n5666)
         );
  OAI22_X1 U2629 ( .A1(n3116), .A2(n3623), .B1(n3314), .B2(n2301), .ZN(n5667)
         );
  OAI22_X1 U2630 ( .A1(n3108), .A2(n3623), .B1(n3314), .B2(n2300), .ZN(n5668)
         );
  OAI22_X1 U2631 ( .A1(n3096), .A2(n3623), .B1(n3314), .B2(n2299), .ZN(n5669)
         );
  OAI22_X1 U2632 ( .A1(n3084), .A2(n3623), .B1(n3314), .B2(n2298), .ZN(n5670)
         );
  OAI22_X1 U2633 ( .A1(n3075), .A2(n3623), .B1(n3314), .B2(n2297), .ZN(n5671)
         );
  OAI22_X1 U2634 ( .A1(n3138), .A2(n3624), .B1(n7134), .B2(n2296), .ZN(n5672)
         );
  OAI22_X1 U2635 ( .A1(n3132), .A2(n3624), .B1(n7134), .B2(n2295), .ZN(n5673)
         );
  OAI22_X1 U2636 ( .A1(n3122), .A2(n3624), .B1(n7134), .B2(n2294), .ZN(n5674)
         );
  OAI22_X1 U2637 ( .A1(n3116), .A2(n3624), .B1(n7134), .B2(n2293), .ZN(n5675)
         );
  OAI22_X1 U2638 ( .A1(n3108), .A2(n3624), .B1(n7134), .B2(n2292), .ZN(n5676)
         );
  OAI22_X1 U2639 ( .A1(n3095), .A2(n3624), .B1(n7134), .B2(n2291), .ZN(n5677)
         );
  OAI22_X1 U2640 ( .A1(n3087), .A2(n3624), .B1(n7134), .B2(n2290), .ZN(n5678)
         );
  OAI22_X1 U2641 ( .A1(n3078), .A2(n3624), .B1(n7134), .B2(n2289), .ZN(n5679)
         );
  OAI22_X1 U2642 ( .A1(n3138), .A2(n3625), .B1(n3234), .B2(n2272), .ZN(n5680)
         );
  OAI22_X1 U2643 ( .A1(n3132), .A2(n3625), .B1(n3234), .B2(n2271), .ZN(n5681)
         );
  OAI22_X1 U2644 ( .A1(n3125), .A2(n3625), .B1(n3234), .B2(n2270), .ZN(n5682)
         );
  OAI22_X1 U2645 ( .A1(n3116), .A2(n3625), .B1(n3234), .B2(n2269), .ZN(n5683)
         );
  OAI22_X1 U2646 ( .A1(n3108), .A2(n3625), .B1(n3234), .B2(n2268), .ZN(n5684)
         );
  OAI22_X1 U2647 ( .A1(n3096), .A2(n3625), .B1(n3234), .B2(n2267), .ZN(n5685)
         );
  OAI22_X1 U2648 ( .A1(n3088), .A2(n3625), .B1(n3234), .B2(n2266), .ZN(n5686)
         );
  OAI22_X1 U2649 ( .A1(n3079), .A2(n3625), .B1(n3234), .B2(n2265), .ZN(n5687)
         );
  OAI22_X1 U2650 ( .A1(n3138), .A2(n3626), .B1(n7182), .B2(n2264), .ZN(n5688)
         );
  OAI22_X1 U2651 ( .A1(n3132), .A2(n3626), .B1(n7182), .B2(n2263), .ZN(n5689)
         );
  OAI22_X1 U2652 ( .A1(n3126), .A2(n3626), .B1(n7182), .B2(n2262), .ZN(n5690)
         );
  OAI22_X1 U2653 ( .A1(n3116), .A2(n3626), .B1(n7182), .B2(n2261), .ZN(n5691)
         );
  OAI22_X1 U2654 ( .A1(n3108), .A2(n3626), .B1(n7182), .B2(n2260), .ZN(n5692)
         );
  OAI22_X1 U2655 ( .A1(n3095), .A2(n3626), .B1(n7182), .B2(n2259), .ZN(n5693)
         );
  OAI22_X1 U2656 ( .A1(n3089), .A2(n3626), .B1(n7182), .B2(n2258), .ZN(n5694)
         );
  OAI22_X1 U2657 ( .A1(n3080), .A2(n3626), .B1(n7182), .B2(n2257), .ZN(n5695)
         );
  OAI22_X1 U2658 ( .A1(n3138), .A2(n3627), .B1(n3298), .B2(n2240), .ZN(n5696)
         );
  OAI22_X1 U2659 ( .A1(n3132), .A2(n3627), .B1(n3298), .B2(n2239), .ZN(n5697)
         );
  OAI22_X1 U2660 ( .A1(n3125), .A2(n3627), .B1(n3298), .B2(n2238), .ZN(n5698)
         );
  OAI22_X1 U2661 ( .A1(n3116), .A2(n3627), .B1(n3298), .B2(n2237), .ZN(n5699)
         );
  OAI22_X1 U2662 ( .A1(n3108), .A2(n3627), .B1(n3298), .B2(n2236), .ZN(n5700)
         );
  OAI22_X1 U2663 ( .A1(n3096), .A2(n3627), .B1(n3298), .B2(n2235), .ZN(n5701)
         );
  OAI22_X1 U2664 ( .A1(n3089), .A2(n3627), .B1(n3298), .B2(n2234), .ZN(n5702)
         );
  OAI22_X1 U2665 ( .A1(n3080), .A2(n3627), .B1(n3298), .B2(n2233), .ZN(n5703)
         );
  OAI22_X1 U2666 ( .A1(n3137), .A2(n3629), .B1(n7118), .B2(n2232), .ZN(n5704)
         );
  OAI22_X1 U2667 ( .A1(n3131), .A2(n3629), .B1(n7118), .B2(n2231), .ZN(n5705)
         );
  OAI22_X1 U2668 ( .A1(n3123), .A2(n3629), .B1(n7118), .B2(n2230), .ZN(n5706)
         );
  OAI22_X1 U2669 ( .A1(n3116), .A2(n3629), .B1(n7118), .B2(n2229), .ZN(n5707)
         );
  OAI22_X1 U2670 ( .A1(n3108), .A2(n3629), .B1(n7118), .B2(n2228), .ZN(n5708)
         );
  OAI22_X1 U2671 ( .A1(n3095), .A2(n3629), .B1(n7118), .B2(n2227), .ZN(n5709)
         );
  OAI22_X1 U2672 ( .A1(n3085), .A2(n3629), .B1(n7118), .B2(n2226), .ZN(n5710)
         );
  OAI22_X1 U2673 ( .A1(n3076), .A2(n3629), .B1(n7118), .B2(n2225), .ZN(n5711)
         );
  OAI22_X1 U2674 ( .A1(n3137), .A2(n3630), .B1(n3281), .B2(n2208), .ZN(n5712)
         );
  OAI22_X1 U2675 ( .A1(n3131), .A2(n3630), .B1(n3281), .B2(n2207), .ZN(n5713)
         );
  OAI22_X1 U2676 ( .A1(n3124), .A2(n3630), .B1(n3281), .B2(n2206), .ZN(n5714)
         );
  OAI22_X1 U2677 ( .A1(n3116), .A2(n3630), .B1(n3281), .B2(n2205), .ZN(n5715)
         );
  OAI22_X1 U2678 ( .A1(n3108), .A2(n3630), .B1(n3281), .B2(n2204), .ZN(n5716)
         );
  OAI22_X1 U2679 ( .A1(n3096), .A2(n3630), .B1(n3281), .B2(n2203), .ZN(n5717)
         );
  OAI22_X1 U2680 ( .A1(n3082), .A2(n3630), .B1(n3281), .B2(n2202), .ZN(n5718)
         );
  OAI22_X1 U2681 ( .A1(n3073), .A2(n3630), .B1(n3281), .B2(n2201), .ZN(n5719)
         );
  OAI22_X1 U2682 ( .A1(n3138), .A2(n3633), .B1(n7229), .B2(n2200), .ZN(n5720)
         );
  OAI22_X1 U2683 ( .A1(n3131), .A2(n3633), .B1(n7229), .B2(n2199), .ZN(n5721)
         );
  OAI22_X1 U2684 ( .A1(n3123), .A2(n3633), .B1(n7229), .B2(n2198), .ZN(n5722)
         );
  OAI22_X1 U2685 ( .A1(n3116), .A2(n3633), .B1(n7229), .B2(n2197), .ZN(n5723)
         );
  OAI22_X1 U2686 ( .A1(n3108), .A2(n3633), .B1(n7229), .B2(n2196), .ZN(n5724)
         );
  OAI22_X1 U2687 ( .A1(n3095), .A2(n3633), .B1(n7229), .B2(n2195), .ZN(n5725)
         );
  OAI22_X1 U2688 ( .A1(n3085), .A2(n3633), .B1(n7229), .B2(n2194), .ZN(n5726)
         );
  OAI22_X1 U2689 ( .A1(n3076), .A2(n3633), .B1(n7229), .B2(n2193), .ZN(n5727)
         );
  OAI22_X1 U2690 ( .A1(n7258), .A2(n3635), .B1(n3345), .B2(n2176), .ZN(n5728)
         );
  OAI22_X1 U2691 ( .A1(n3131), .A2(n3635), .B1(n3345), .B2(n2175), .ZN(n5729)
         );
  OAI22_X1 U2692 ( .A1(n3124), .A2(n3635), .B1(n3345), .B2(n2174), .ZN(n5730)
         );
  OAI22_X1 U2693 ( .A1(n3116), .A2(n3635), .B1(n3345), .B2(n2173), .ZN(n5731)
         );
  OAI22_X1 U2694 ( .A1(n3108), .A2(n3635), .B1(n3345), .B2(n2172), .ZN(n5732)
         );
  OAI22_X1 U2695 ( .A1(n3096), .A2(n3635), .B1(n3345), .B2(n2171), .ZN(n5733)
         );
  OAI22_X1 U2696 ( .A1(n3086), .A2(n3635), .B1(n3345), .B2(n2170), .ZN(n5734)
         );
  OAI22_X1 U2697 ( .A1(n3077), .A2(n3635), .B1(n3345), .B2(n2169), .ZN(n5735)
         );
  OAI22_X1 U2698 ( .A1(n3138), .A2(n3638), .B1(n7165), .B2(n2168), .ZN(n5736)
         );
  OAI22_X1 U2699 ( .A1(n3131), .A2(n3638), .B1(n7165), .B2(n2167), .ZN(n5737)
         );
  OAI22_X1 U2700 ( .A1(n3123), .A2(n3638), .B1(n7165), .B2(n2166), .ZN(n5738)
         );
  OAI22_X1 U2701 ( .A1(n3116), .A2(n3638), .B1(n7165), .B2(n2165), .ZN(n5739)
         );
  OAI22_X1 U2702 ( .A1(n3108), .A2(n3638), .B1(n7165), .B2(n2164), .ZN(n5740)
         );
  OAI22_X1 U2703 ( .A1(n3097), .A2(n3638), .B1(n7165), .B2(n2163), .ZN(n5741)
         );
  OAI22_X1 U2704 ( .A1(n3082), .A2(n3638), .B1(n7165), .B2(n2162), .ZN(n5742)
         );
  OAI22_X1 U2705 ( .A1(n3073), .A2(n3638), .B1(n7165), .B2(n2161), .ZN(n5743)
         );
  OAI22_X1 U2706 ( .A1(n3138), .A2(n3640), .B1(n3265), .B2(n2144), .ZN(n5744)
         );
  OAI22_X1 U2707 ( .A1(n3131), .A2(n3640), .B1(n3265), .B2(n2143), .ZN(n5745)
         );
  OAI22_X1 U2708 ( .A1(n3124), .A2(n3640), .B1(n3265), .B2(n2142), .ZN(n5746)
         );
  OAI22_X1 U2709 ( .A1(n3116), .A2(n3640), .B1(n3265), .B2(n2141), .ZN(n5747)
         );
  OAI22_X1 U2710 ( .A1(n3108), .A2(n3640), .B1(n3265), .B2(n2140), .ZN(n5748)
         );
  OAI22_X1 U2711 ( .A1(n3091), .A2(n3640), .B1(n3265), .B2(n2139), .ZN(n5749)
         );
  OAI22_X1 U2712 ( .A1(n3089), .A2(n3640), .B1(n3265), .B2(n2138), .ZN(n5750)
         );
  OAI22_X1 U2713 ( .A1(n3080), .A2(n3640), .B1(n3265), .B2(n2137), .ZN(n5751)
         );
  OAI22_X1 U2714 ( .A1(n3137), .A2(n3641), .B1(n7213), .B2(n2136), .ZN(n5752)
         );
  OAI22_X1 U2715 ( .A1(n3131), .A2(n3641), .B1(n7213), .B2(n2135), .ZN(n5753)
         );
  OAI22_X1 U2716 ( .A1(n3123), .A2(n3641), .B1(n7213), .B2(n2134), .ZN(n5754)
         );
  OAI22_X1 U2717 ( .A1(n3116), .A2(n3641), .B1(n7213), .B2(n2133), .ZN(n5755)
         );
  OAI22_X1 U2718 ( .A1(n3108), .A2(n3641), .B1(n7213), .B2(n2132), .ZN(n5756)
         );
  OAI22_X1 U2719 ( .A1(n3095), .A2(n3641), .B1(n7213), .B2(n2131), .ZN(n5757)
         );
  OAI22_X1 U2720 ( .A1(n3090), .A2(n3641), .B1(n7213), .B2(n2130), .ZN(n5758)
         );
  OAI22_X1 U2721 ( .A1(n3081), .A2(n3641), .B1(n7213), .B2(n2129), .ZN(n5759)
         );
  OAI22_X1 U2722 ( .A1(n3144), .A2(n3642), .B1(n3329), .B2(n2112), .ZN(n5760)
         );
  OAI22_X1 U2723 ( .A1(n3131), .A2(n3642), .B1(n3329), .B2(n2111), .ZN(n5761)
         );
  OAI22_X1 U2724 ( .A1(n3124), .A2(n3642), .B1(n3329), .B2(n2110), .ZN(n5762)
         );
  OAI22_X1 U2725 ( .A1(n3117), .A2(n3642), .B1(n3329), .B2(n2109), .ZN(n5763)
         );
  OAI22_X1 U2726 ( .A1(n3105), .A2(n3642), .B1(n3329), .B2(n2108), .ZN(n5764)
         );
  OAI22_X1 U2727 ( .A1(n3094), .A2(n3642), .B1(n3329), .B2(n2107), .ZN(n5765)
         );
  OAI22_X1 U2728 ( .A1(n3090), .A2(n3642), .B1(n3329), .B2(n2106), .ZN(n5766)
         );
  OAI22_X1 U2729 ( .A1(n3081), .A2(n3642), .B1(n3329), .B2(n2105), .ZN(n5767)
         );
  OAI22_X1 U2730 ( .A1(n3143), .A2(n3644), .B1(n7149), .B2(n2104), .ZN(n5768)
         );
  OAI22_X1 U2731 ( .A1(n3131), .A2(n3644), .B1(n7149), .B2(n2103), .ZN(n5769)
         );
  OAI22_X1 U2732 ( .A1(n3123), .A2(n3644), .B1(n7149), .B2(n2102), .ZN(n5770)
         );
  OAI22_X1 U2733 ( .A1(n3117), .A2(n3644), .B1(n7149), .B2(n2101), .ZN(n5771)
         );
  OAI22_X1 U2734 ( .A1(n3101), .A2(n3644), .B1(n7149), .B2(n2100), .ZN(n5772)
         );
  OAI22_X1 U2735 ( .A1(n3094), .A2(n3644), .B1(n7149), .B2(n2099), .ZN(n5773)
         );
  OAI22_X1 U2736 ( .A1(n3090), .A2(n3644), .B1(n7149), .B2(n2098), .ZN(n5774)
         );
  OAI22_X1 U2737 ( .A1(n3081), .A2(n3644), .B1(n7149), .B2(n2097), .ZN(n5775)
         );
  OAI22_X1 U2738 ( .A1(n3142), .A2(n3645), .B1(n3249), .B2(n2080), .ZN(n5776)
         );
  OAI22_X1 U2739 ( .A1(n3131), .A2(n3645), .B1(n3249), .B2(n2079), .ZN(n5777)
         );
  OAI22_X1 U2740 ( .A1(n3124), .A2(n3645), .B1(n3249), .B2(n2078), .ZN(n5778)
         );
  OAI22_X1 U2741 ( .A1(n3117), .A2(n3645), .B1(n3249), .B2(n2077), .ZN(n5779)
         );
  OAI22_X1 U2742 ( .A1(n3105), .A2(n3645), .B1(n3249), .B2(n2076), .ZN(n5780)
         );
  OAI22_X1 U2743 ( .A1(n3094), .A2(n3645), .B1(n3249), .B2(n2075), .ZN(n5781)
         );
  OAI22_X1 U2744 ( .A1(n3090), .A2(n3645), .B1(n3249), .B2(n2074), .ZN(n5782)
         );
  OAI22_X1 U2745 ( .A1(n3081), .A2(n3645), .B1(n3249), .B2(n2073), .ZN(n5783)
         );
  OAI22_X1 U2746 ( .A1(n3145), .A2(n3646), .B1(n7197), .B2(n2072), .ZN(n5784)
         );
  OAI22_X1 U2747 ( .A1(n3131), .A2(n3646), .B1(n7197), .B2(n2071), .ZN(n5785)
         );
  OAI22_X1 U2748 ( .A1(n3123), .A2(n3646), .B1(n7197), .B2(n2070), .ZN(n5786)
         );
  OAI22_X1 U2749 ( .A1(n3117), .A2(n3646), .B1(n7197), .B2(n2069), .ZN(n5787)
         );
  OAI22_X1 U2750 ( .A1(n3104), .A2(n3646), .B1(n7197), .B2(n2068), .ZN(n5788)
         );
  OAI22_X1 U2751 ( .A1(n3094), .A2(n3646), .B1(n7197), .B2(n2067), .ZN(n5789)
         );
  OAI22_X1 U2752 ( .A1(n3090), .A2(n3646), .B1(n7197), .B2(n2066), .ZN(n5790)
         );
  OAI22_X1 U2753 ( .A1(n3081), .A2(n3646), .B1(n7197), .B2(n2065), .ZN(n5791)
         );
  OAI22_X1 U2754 ( .A1(n3144), .A2(n3647), .B1(n3313), .B2(n2048), .ZN(n5792)
         );
  OAI22_X1 U2755 ( .A1(n3131), .A2(n3647), .B1(n3313), .B2(n2047), .ZN(n5793)
         );
  OAI22_X1 U2756 ( .A1(n3124), .A2(n3647), .B1(n3313), .B2(n2046), .ZN(n5794)
         );
  OAI22_X1 U2757 ( .A1(n3117), .A2(n3647), .B1(n3313), .B2(n2045), .ZN(n5795)
         );
  OAI22_X1 U2758 ( .A1(n3105), .A2(n3647), .B1(n3313), .B2(n2044), .ZN(n5796)
         );
  OAI22_X1 U2759 ( .A1(n3097), .A2(n3647), .B1(n3313), .B2(n2043), .ZN(n5797)
         );
  OAI22_X1 U2760 ( .A1(n3090), .A2(n3647), .B1(n3313), .B2(n2042), .ZN(n5798)
         );
  OAI22_X1 U2761 ( .A1(n3081), .A2(n3647), .B1(n3313), .B2(n2041), .ZN(n5799)
         );
  OAI22_X1 U2762 ( .A1(n3143), .A2(n3649), .B1(n7133), .B2(n2040), .ZN(n5800)
         );
  OAI22_X1 U2763 ( .A1(n3131), .A2(n3649), .B1(n7133), .B2(n2039), .ZN(n5801)
         );
  OAI22_X1 U2764 ( .A1(n3126), .A2(n3649), .B1(n7133), .B2(n2038), .ZN(n5802)
         );
  OAI22_X1 U2765 ( .A1(n3117), .A2(n3649), .B1(n7133), .B2(n2037), .ZN(n5803)
         );
  OAI22_X1 U2766 ( .A1(n3101), .A2(n3649), .B1(n7133), .B2(n2036), .ZN(n5804)
         );
  OAI22_X1 U2767 ( .A1(n3097), .A2(n3649), .B1(n7133), .B2(n2035), .ZN(n5805)
         );
  OAI22_X1 U2768 ( .A1(n3090), .A2(n3649), .B1(n7133), .B2(n2034), .ZN(n5806)
         );
  OAI22_X1 U2769 ( .A1(n3081), .A2(n3649), .B1(n7133), .B2(n2033), .ZN(n5807)
         );
  OAI22_X1 U2770 ( .A1(n3139), .A2(n3650), .B1(n3233), .B2(n2016), .ZN(n5808)
         );
  OAI22_X1 U2771 ( .A1(n3134), .A2(n3650), .B1(n3233), .B2(n2015), .ZN(n5809)
         );
  OAI22_X1 U2772 ( .A1(n3120), .A2(n3650), .B1(n3233), .B2(n2014), .ZN(n5810)
         );
  OAI22_X1 U2773 ( .A1(n3117), .A2(n3650), .B1(n3233), .B2(n2013), .ZN(n5811)
         );
  OAI22_X1 U2774 ( .A1(n3104), .A2(n3650), .B1(n3233), .B2(n2012), .ZN(n5812)
         );
  OAI22_X1 U2775 ( .A1(n3097), .A2(n3650), .B1(n3233), .B2(n2011), .ZN(n5813)
         );
  OAI22_X1 U2776 ( .A1(n3090), .A2(n3650), .B1(n3233), .B2(n2010), .ZN(n5814)
         );
  OAI22_X1 U2777 ( .A1(n3081), .A2(n3650), .B1(n3233), .B2(n2009), .ZN(n5815)
         );
  OAI22_X1 U2778 ( .A1(n3140), .A2(n3651), .B1(n7181), .B2(n2008), .ZN(n5816)
         );
  OAI22_X1 U2779 ( .A1(n3131), .A2(n3651), .B1(n7181), .B2(n2007), .ZN(n5817)
         );
  OAI22_X1 U2780 ( .A1(n3123), .A2(n3651), .B1(n7181), .B2(n2006), .ZN(n5818)
         );
  OAI22_X1 U2781 ( .A1(n3117), .A2(n3651), .B1(n7181), .B2(n2005), .ZN(n5819)
         );
  OAI22_X1 U2782 ( .A1(n3101), .A2(n3651), .B1(n7181), .B2(n2004), .ZN(n5820)
         );
  OAI22_X1 U2783 ( .A1(n3097), .A2(n3651), .B1(n7181), .B2(n2003), .ZN(n5821)
         );
  OAI22_X1 U2784 ( .A1(n3090), .A2(n3651), .B1(n7181), .B2(n2002), .ZN(n5822)
         );
  OAI22_X1 U2785 ( .A1(n3081), .A2(n3651), .B1(n7181), .B2(n2001), .ZN(n5823)
         );
  OAI22_X1 U2786 ( .A1(n7258), .A2(n3382), .B1(n7132), .B2(n1720), .ZN(n5960)
         );
  OAI22_X1 U2787 ( .A1(n3129), .A2(n3382), .B1(n7132), .B2(n1719), .ZN(n5961)
         );
  OAI22_X1 U2788 ( .A1(n3119), .A2(n3382), .B1(n7132), .B2(n1718), .ZN(n5962)
         );
  OAI22_X1 U2789 ( .A1(n3116), .A2(n3382), .B1(n7132), .B2(n1717), .ZN(n5963)
         );
  OAI22_X1 U2790 ( .A1(n3106), .A2(n3382), .B1(n7132), .B2(n1716), .ZN(n5964)
         );
  OAI22_X1 U2791 ( .A1(n3091), .A2(n3382), .B1(n7132), .B2(n1715), .ZN(n5965)
         );
  OAI22_X1 U2792 ( .A1(n3082), .A2(n3382), .B1(n7132), .B2(n1714), .ZN(n5966)
         );
  OAI22_X1 U2793 ( .A1(n3073), .A2(n3382), .B1(n7132), .B2(n1713), .ZN(n5967)
         );
  OAI22_X1 U2794 ( .A1(n7258), .A2(n3384), .B1(n3295), .B2(n1696), .ZN(n5968)
         );
  OAI22_X1 U2795 ( .A1(n3132), .A2(n3384), .B1(n3295), .B2(n1695), .ZN(n5969)
         );
  OAI22_X1 U2796 ( .A1(n3120), .A2(n3384), .B1(n3295), .B2(n1694), .ZN(n5970)
         );
  OAI22_X1 U2797 ( .A1(n7255), .A2(n3384), .B1(n3295), .B2(n1693), .ZN(n5971)
         );
  OAI22_X1 U2798 ( .A1(n7254), .A2(n3384), .B1(n3295), .B2(n1692), .ZN(n5972)
         );
  OAI22_X1 U2799 ( .A1(n3093), .A2(n3384), .B1(n3295), .B2(n1691), .ZN(n5973)
         );
  OAI22_X1 U2800 ( .A1(n3082), .A2(n3384), .B1(n3295), .B2(n1690), .ZN(n5974)
         );
  OAI22_X1 U2801 ( .A1(n3073), .A2(n3384), .B1(n3295), .B2(n1689), .ZN(n5975)
         );
  OAI22_X1 U2802 ( .A1(n7258), .A2(n3385), .B1(n7243), .B2(n1688), .ZN(n5976)
         );
  OAI22_X1 U2803 ( .A1(n3130), .A2(n3385), .B1(n7243), .B2(n1687), .ZN(n5977)
         );
  OAI22_X1 U2804 ( .A1(n3118), .A2(n3385), .B1(n7243), .B2(n1686), .ZN(n5978)
         );
  OAI22_X1 U2805 ( .A1(n7255), .A2(n3385), .B1(n7243), .B2(n1685), .ZN(n5979)
         );
  OAI22_X1 U2806 ( .A1(n7254), .A2(n3385), .B1(n7243), .B2(n1684), .ZN(n5980)
         );
  OAI22_X1 U2807 ( .A1(n3096), .A2(n3385), .B1(n7243), .B2(n1683), .ZN(n5981)
         );
  OAI22_X1 U2808 ( .A1(n3083), .A2(n3385), .B1(n7243), .B2(n1682), .ZN(n5982)
         );
  OAI22_X1 U2809 ( .A1(n3074), .A2(n3385), .B1(n7243), .B2(n1681), .ZN(n5983)
         );
  OAI22_X1 U2810 ( .A1(n7258), .A2(n3386), .B1(n7114), .B2(n1664), .ZN(n5984)
         );
  OAI22_X1 U2811 ( .A1(n7257), .A2(n3386), .B1(n7114), .B2(n1663), .ZN(n5985)
         );
  OAI22_X1 U2812 ( .A1(n3118), .A2(n3386), .B1(n7114), .B2(n1662), .ZN(n5986)
         );
  OAI22_X1 U2813 ( .A1(n7255), .A2(n3386), .B1(n7114), .B2(n1661), .ZN(n5987)
         );
  OAI22_X1 U2814 ( .A1(n7254), .A2(n3386), .B1(n7114), .B2(n1660), .ZN(n5988)
         );
  OAI22_X1 U2815 ( .A1(n7253), .A2(n3386), .B1(n7114), .B2(n1659), .ZN(n5989)
         );
  OAI22_X1 U2816 ( .A1(n7252), .A2(n3386), .B1(n7114), .B2(n1658), .ZN(n5990)
         );
  OAI22_X1 U2817 ( .A1(n7251), .A2(n3386), .B1(n7114), .B2(n1657), .ZN(n5991)
         );
  OAI22_X1 U2818 ( .A1(n7258), .A2(n3387), .B1(n7179), .B2(n1656), .ZN(n5992)
         );
  OAI22_X1 U2819 ( .A1(n7257), .A2(n3387), .B1(n7179), .B2(n1655), .ZN(n5993)
         );
  OAI22_X1 U2820 ( .A1(n3118), .A2(n3387), .B1(n7179), .B2(n1654), .ZN(n5994)
         );
  OAI22_X1 U2821 ( .A1(n7255), .A2(n3387), .B1(n7179), .B2(n1653), .ZN(n5995)
         );
  OAI22_X1 U2822 ( .A1(n7254), .A2(n3387), .B1(n7179), .B2(n1652), .ZN(n5996)
         );
  OAI22_X1 U2823 ( .A1(n3091), .A2(n3387), .B1(n7179), .B2(n1651), .ZN(n5997)
         );
  OAI22_X1 U2824 ( .A1(n3083), .A2(n3387), .B1(n7179), .B2(n1650), .ZN(n5998)
         );
  OAI22_X1 U2825 ( .A1(n3074), .A2(n3387), .B1(n7179), .B2(n1649), .ZN(n5999)
         );
  OAI22_X1 U2826 ( .A1(n7258), .A2(n3388), .B1(n3279), .B2(n1632), .ZN(n6000)
         );
  OAI22_X1 U2827 ( .A1(n7257), .A2(n3388), .B1(n3279), .B2(n1631), .ZN(n6001)
         );
  OAI22_X1 U2828 ( .A1(n3118), .A2(n3388), .B1(n3279), .B2(n1630), .ZN(n6002)
         );
  OAI22_X1 U2829 ( .A1(n7255), .A2(n3388), .B1(n3279), .B2(n1629), .ZN(n6003)
         );
  OAI22_X1 U2830 ( .A1(n7254), .A2(n3388), .B1(n3279), .B2(n1628), .ZN(n6004)
         );
  OAI22_X1 U2831 ( .A1(n3099), .A2(n3388), .B1(n3279), .B2(n1627), .ZN(n6005)
         );
  OAI22_X1 U2832 ( .A1(n3087), .A2(n3388), .B1(n3279), .B2(n1626), .ZN(n6006)
         );
  OAI22_X1 U2833 ( .A1(n3078), .A2(n3388), .B1(n3279), .B2(n1625), .ZN(n6007)
         );
  OAI22_X1 U2834 ( .A1(n7258), .A2(n3389), .B1(n7227), .B2(n1624), .ZN(n6008)
         );
  OAI22_X1 U2835 ( .A1(n7257), .A2(n3389), .B1(n7227), .B2(n1623), .ZN(n6009)
         );
  OAI22_X1 U2836 ( .A1(n3119), .A2(n3389), .B1(n7227), .B2(n1622), .ZN(n6010)
         );
  OAI22_X1 U2837 ( .A1(n7255), .A2(n3389), .B1(n7227), .B2(n1621), .ZN(n6011)
         );
  OAI22_X1 U2838 ( .A1(n7254), .A2(n3389), .B1(n7227), .B2(n1620), .ZN(n6012)
         );
  OAI22_X1 U2839 ( .A1(n3091), .A2(n3389), .B1(n7227), .B2(n1619), .ZN(n6013)
         );
  OAI22_X1 U2840 ( .A1(n7252), .A2(n3389), .B1(n7227), .B2(n1618), .ZN(n6014)
         );
  OAI22_X1 U2841 ( .A1(n7251), .A2(n3389), .B1(n7227), .B2(n1617), .ZN(n6015)
         );
  OAI22_X1 U2842 ( .A1(n7258), .A2(n3390), .B1(n3343), .B2(n1600), .ZN(n6016)
         );
  OAI22_X1 U2843 ( .A1(n7257), .A2(n3390), .B1(n3343), .B2(n1599), .ZN(n6017)
         );
  OAI22_X1 U2844 ( .A1(n3119), .A2(n3390), .B1(n3343), .B2(n1598), .ZN(n6018)
         );
  OAI22_X1 U2845 ( .A1(n7255), .A2(n3390), .B1(n3343), .B2(n1597), .ZN(n6019)
         );
  OAI22_X1 U2846 ( .A1(n7254), .A2(n3390), .B1(n3343), .B2(n1596), .ZN(n6020)
         );
  OAI22_X1 U2847 ( .A1(n3093), .A2(n3390), .B1(n3343), .B2(n1595), .ZN(n6021)
         );
  OAI22_X1 U2848 ( .A1(n7252), .A2(n3390), .B1(n3343), .B2(n1594), .ZN(n6022)
         );
  OAI22_X1 U2849 ( .A1(n7251), .A2(n3390), .B1(n3343), .B2(n1593), .ZN(n6023)
         );
  OAI22_X1 U2850 ( .A1(n7258), .A2(n3391), .B1(n7163), .B2(n1592), .ZN(n6024)
         );
  OAI22_X1 U2851 ( .A1(n7257), .A2(n3391), .B1(n7163), .B2(n1591), .ZN(n6025)
         );
  OAI22_X1 U2852 ( .A1(n3119), .A2(n3391), .B1(n7163), .B2(n1590), .ZN(n6026)
         );
  OAI22_X1 U2853 ( .A1(n7255), .A2(n3391), .B1(n7163), .B2(n1589), .ZN(n6027)
         );
  OAI22_X1 U2854 ( .A1(n7254), .A2(n3391), .B1(n7163), .B2(n1588), .ZN(n6028)
         );
  OAI22_X1 U2855 ( .A1(n3098), .A2(n3391), .B1(n7163), .B2(n1587), .ZN(n6029)
         );
  OAI22_X1 U2856 ( .A1(n7252), .A2(n3391), .B1(n7163), .B2(n1586), .ZN(n6030)
         );
  OAI22_X1 U2857 ( .A1(n7251), .A2(n3391), .B1(n7163), .B2(n1585), .ZN(n6031)
         );
  OAI22_X1 U2858 ( .A1(n7258), .A2(n3392), .B1(n3263), .B2(n1568), .ZN(n6032)
         );
  OAI22_X1 U2859 ( .A1(n7257), .A2(n3392), .B1(n3263), .B2(n1567), .ZN(n6033)
         );
  OAI22_X1 U2860 ( .A1(n3119), .A2(n3392), .B1(n3263), .B2(n1566), .ZN(n6034)
         );
  OAI22_X1 U2861 ( .A1(n7255), .A2(n3392), .B1(n3263), .B2(n1565), .ZN(n6035)
         );
  OAI22_X1 U2862 ( .A1(n7254), .A2(n3392), .B1(n3263), .B2(n1564), .ZN(n6036)
         );
  OAI22_X1 U2863 ( .A1(n3091), .A2(n3392), .B1(n3263), .B2(n1563), .ZN(n6037)
         );
  OAI22_X1 U2864 ( .A1(n7252), .A2(n3392), .B1(n3263), .B2(n1562), .ZN(n6038)
         );
  OAI22_X1 U2865 ( .A1(n7251), .A2(n3392), .B1(n3263), .B2(n1561), .ZN(n6039)
         );
  OAI22_X1 U2866 ( .A1(n7258), .A2(n3393), .B1(n7211), .B2(n1560), .ZN(n6040)
         );
  OAI22_X1 U2867 ( .A1(n3136), .A2(n3393), .B1(n7211), .B2(n1559), .ZN(n6041)
         );
  OAI22_X1 U2868 ( .A1(n3120), .A2(n3393), .B1(n7211), .B2(n1558), .ZN(n6042)
         );
  OAI22_X1 U2869 ( .A1(n3110), .A2(n3393), .B1(n7211), .B2(n1557), .ZN(n6043)
         );
  OAI22_X1 U2870 ( .A1(n3105), .A2(n3393), .B1(n7211), .B2(n1556), .ZN(n6044)
         );
  OAI22_X1 U2871 ( .A1(n3093), .A2(n3393), .B1(n7211), .B2(n1555), .ZN(n6045)
         );
  OAI22_X1 U2872 ( .A1(n3083), .A2(n3393), .B1(n7211), .B2(n1554), .ZN(n6046)
         );
  OAI22_X1 U2873 ( .A1(n3074), .A2(n3393), .B1(n7211), .B2(n1553), .ZN(n6047)
         );
  OAI22_X1 U2874 ( .A1(n7258), .A2(n3394), .B1(n3327), .B2(n1536), .ZN(n6048)
         );
  OAI22_X1 U2875 ( .A1(n3136), .A2(n3394), .B1(n3327), .B2(n1535), .ZN(n6049)
         );
  OAI22_X1 U2876 ( .A1(n3119), .A2(n3394), .B1(n3327), .B2(n1534), .ZN(n6050)
         );
  OAI22_X1 U2877 ( .A1(n7255), .A2(n3394), .B1(n3327), .B2(n1533), .ZN(n6051)
         );
  OAI22_X1 U2878 ( .A1(n3105), .A2(n3394), .B1(n3327), .B2(n1532), .ZN(n6052)
         );
  OAI22_X1 U2879 ( .A1(n3099), .A2(n3394), .B1(n3327), .B2(n1531), .ZN(n6053)
         );
  OAI22_X1 U2880 ( .A1(n7252), .A2(n3394), .B1(n3327), .B2(n1530), .ZN(n6054)
         );
  OAI22_X1 U2881 ( .A1(n7251), .A2(n3394), .B1(n3327), .B2(n1529), .ZN(n6055)
         );
  OAI22_X1 U2882 ( .A1(n3144), .A2(n3395), .B1(n7147), .B2(n1528), .ZN(n6056)
         );
  OAI22_X1 U2883 ( .A1(n3136), .A2(n3395), .B1(n7147), .B2(n1527), .ZN(n6057)
         );
  OAI22_X1 U2884 ( .A1(n3118), .A2(n3395), .B1(n7147), .B2(n1526), .ZN(n6058)
         );
  OAI22_X1 U2885 ( .A1(n3110), .A2(n3395), .B1(n7147), .B2(n1525), .ZN(n6059)
         );
  OAI22_X1 U2886 ( .A1(n3105), .A2(n3395), .B1(n7147), .B2(n1524), .ZN(n6060)
         );
  OAI22_X1 U2887 ( .A1(n3093), .A2(n3395), .B1(n7147), .B2(n1523), .ZN(n6061)
         );
  OAI22_X1 U2888 ( .A1(n3088), .A2(n3395), .B1(n7147), .B2(n1522), .ZN(n6062)
         );
  OAI22_X1 U2889 ( .A1(n3079), .A2(n3395), .B1(n7147), .B2(n1521), .ZN(n6063)
         );
  OAI22_X1 U2890 ( .A1(n3143), .A2(n3396), .B1(n3247), .B2(n1504), .ZN(n6064)
         );
  OAI22_X1 U2891 ( .A1(n3128), .A2(n3396), .B1(n3247), .B2(n1503), .ZN(n6065)
         );
  OAI22_X1 U2892 ( .A1(n3118), .A2(n3396), .B1(n3247), .B2(n1502), .ZN(n6066)
         );
  OAI22_X1 U2893 ( .A1(n7255), .A2(n3396), .B1(n3247), .B2(n1501), .ZN(n6067)
         );
  OAI22_X1 U2894 ( .A1(n3105), .A2(n3396), .B1(n3247), .B2(n1500), .ZN(n6068)
         );
  OAI22_X1 U2895 ( .A1(n3093), .A2(n3396), .B1(n3247), .B2(n1499), .ZN(n6069)
         );
  OAI22_X1 U2896 ( .A1(n3083), .A2(n3396), .B1(n3247), .B2(n1498), .ZN(n6070)
         );
  OAI22_X1 U2897 ( .A1(n3074), .A2(n3396), .B1(n3247), .B2(n1497), .ZN(n6071)
         );
  OAI22_X1 U2898 ( .A1(n3142), .A2(n3397), .B1(n7195), .B2(n1496), .ZN(n6072)
         );
  OAI22_X1 U2899 ( .A1(n3136), .A2(n3397), .B1(n7195), .B2(n1495), .ZN(n6073)
         );
  OAI22_X1 U2900 ( .A1(n3119), .A2(n3397), .B1(n7195), .B2(n1494), .ZN(n6074)
         );
  OAI22_X1 U2901 ( .A1(n3117), .A2(n3397), .B1(n7195), .B2(n1493), .ZN(n6075)
         );
  OAI22_X1 U2902 ( .A1(n7254), .A2(n3397), .B1(n7195), .B2(n1492), .ZN(n6076)
         );
  OAI22_X1 U2903 ( .A1(n3091), .A2(n3397), .B1(n7195), .B2(n1491), .ZN(n6077)
         );
  OAI22_X1 U2904 ( .A1(n3083), .A2(n3397), .B1(n7195), .B2(n1490), .ZN(n6078)
         );
  OAI22_X1 U2905 ( .A1(n3074), .A2(n3397), .B1(n7195), .B2(n1489), .ZN(n6079)
         );
  OAI22_X1 U2906 ( .A1(n3141), .A2(n3400), .B1(n3311), .B2(n1472), .ZN(n6080)
         );
  OAI22_X1 U2907 ( .A1(n3128), .A2(n3400), .B1(n3311), .B2(n1471), .ZN(n6081)
         );
  OAI22_X1 U2908 ( .A1(n3119), .A2(n3400), .B1(n3311), .B2(n1470), .ZN(n6082)
         );
  OAI22_X1 U2909 ( .A1(n3116), .A2(n3400), .B1(n3311), .B2(n1469), .ZN(n6083)
         );
  OAI22_X1 U2910 ( .A1(n3106), .A2(n3400), .B1(n3311), .B2(n1468), .ZN(n6084)
         );
  OAI22_X1 U2911 ( .A1(n3093), .A2(n3400), .B1(n3311), .B2(n1467), .ZN(n6085)
         );
  OAI22_X1 U2912 ( .A1(n3089), .A2(n3400), .B1(n3311), .B2(n1466), .ZN(n6086)
         );
  OAI22_X1 U2913 ( .A1(n3080), .A2(n3400), .B1(n3311), .B2(n1465), .ZN(n6087)
         );
  OAI22_X1 U2914 ( .A1(n3144), .A2(n3402), .B1(n7131), .B2(n1464), .ZN(n6088)
         );
  OAI22_X1 U2915 ( .A1(n3129), .A2(n3402), .B1(n7131), .B2(n1463), .ZN(n6089)
         );
  OAI22_X1 U2916 ( .A1(n3119), .A2(n3402), .B1(n7131), .B2(n1462), .ZN(n6090)
         );
  OAI22_X1 U2917 ( .A1(n3111), .A2(n3402), .B1(n7131), .B2(n1461), .ZN(n6091)
         );
  OAI22_X1 U2918 ( .A1(n3101), .A2(n3402), .B1(n7131), .B2(n1460), .ZN(n6092)
         );
  OAI22_X1 U2919 ( .A1(n3099), .A2(n3402), .B1(n7131), .B2(n1459), .ZN(n6093)
         );
  OAI22_X1 U2920 ( .A1(n7252), .A2(n3402), .B1(n7131), .B2(n1458), .ZN(n6094)
         );
  OAI22_X1 U2921 ( .A1(n7251), .A2(n3402), .B1(n7131), .B2(n1457), .ZN(n6095)
         );
  OAI22_X1 U2922 ( .A1(n3143), .A2(n3403), .B1(n3294), .B2(n1440), .ZN(n6096)
         );
  OAI22_X1 U2923 ( .A1(n3128), .A2(n3403), .B1(n3294), .B2(n1439), .ZN(n6097)
         );
  OAI22_X1 U2924 ( .A1(n3119), .A2(n3403), .B1(n3294), .B2(n1438), .ZN(n6098)
         );
  OAI22_X1 U2925 ( .A1(n3117), .A2(n3403), .B1(n3294), .B2(n1437), .ZN(n6099)
         );
  OAI22_X1 U2926 ( .A1(n3103), .A2(n3403), .B1(n3294), .B2(n1436), .ZN(n6100)
         );
  OAI22_X1 U2927 ( .A1(n3098), .A2(n3403), .B1(n3294), .B2(n1435), .ZN(n6101)
         );
  OAI22_X1 U2928 ( .A1(n7252), .A2(n3403), .B1(n3294), .B2(n1434), .ZN(n6102)
         );
  OAI22_X1 U2929 ( .A1(n7251), .A2(n3403), .B1(n3294), .B2(n1433), .ZN(n6103)
         );
  OAI22_X1 U2930 ( .A1(n7258), .A2(n3404), .B1(n7242), .B2(n1432), .ZN(n6104)
         );
  OAI22_X1 U2931 ( .A1(n3130), .A2(n3404), .B1(n7242), .B2(n1431), .ZN(n6105)
         );
  OAI22_X1 U2932 ( .A1(n3119), .A2(n3404), .B1(n7242), .B2(n1430), .ZN(n6106)
         );
  OAI22_X1 U2933 ( .A1(n3117), .A2(n3404), .B1(n7242), .B2(n1429), .ZN(n6107)
         );
  OAI22_X1 U2934 ( .A1(n3106), .A2(n3404), .B1(n7242), .B2(n1428), .ZN(n6108)
         );
  OAI22_X1 U2935 ( .A1(n3093), .A2(n3404), .B1(n7242), .B2(n1427), .ZN(n6109)
         );
  OAI22_X1 U2936 ( .A1(n7252), .A2(n3404), .B1(n7242), .B2(n1426), .ZN(n6110)
         );
  OAI22_X1 U2937 ( .A1(n7251), .A2(n3404), .B1(n7242), .B2(n1425), .ZN(n6111)
         );
  OAI22_X1 U2938 ( .A1(n7258), .A2(n3405), .B1(n7113), .B2(n1408), .ZN(n6112)
         );
  OAI22_X1 U2939 ( .A1(n3129), .A2(n3405), .B1(n7113), .B2(n1407), .ZN(n6113)
         );
  OAI22_X1 U2940 ( .A1(n3119), .A2(n3405), .B1(n7113), .B2(n1406), .ZN(n6114)
         );
  OAI22_X1 U2941 ( .A1(n3111), .A2(n3405), .B1(n7113), .B2(n1405), .ZN(n6115)
         );
  OAI22_X1 U2942 ( .A1(n3100), .A2(n3405), .B1(n7113), .B2(n1404), .ZN(n6116)
         );
  OAI22_X1 U2943 ( .A1(n3093), .A2(n3405), .B1(n7113), .B2(n1403), .ZN(n6117)
         );
  OAI22_X1 U2944 ( .A1(n7252), .A2(n3405), .B1(n7113), .B2(n1402), .ZN(n6118)
         );
  OAI22_X1 U2945 ( .A1(n7251), .A2(n3405), .B1(n7113), .B2(n1401), .ZN(n6119)
         );
  OAI22_X1 U2946 ( .A1(n7258), .A2(n3406), .B1(n7178), .B2(n1400), .ZN(n6120)
         );
  OAI22_X1 U2947 ( .A1(n3128), .A2(n3406), .B1(n7178), .B2(n1399), .ZN(n6121)
         );
  OAI22_X1 U2948 ( .A1(n3119), .A2(n3406), .B1(n7178), .B2(n1398), .ZN(n6122)
         );
  OAI22_X1 U2949 ( .A1(n3114), .A2(n3406), .B1(n7178), .B2(n1397), .ZN(n6123)
         );
  OAI22_X1 U2950 ( .A1(n7254), .A2(n3406), .B1(n7178), .B2(n1396), .ZN(n6124)
         );
  OAI22_X1 U2951 ( .A1(n3091), .A2(n3406), .B1(n7178), .B2(n1395), .ZN(n6125)
         );
  OAI22_X1 U2952 ( .A1(n7252), .A2(n3406), .B1(n7178), .B2(n1394), .ZN(n6126)
         );
  OAI22_X1 U2953 ( .A1(n7251), .A2(n3406), .B1(n7178), .B2(n1393), .ZN(n6127)
         );
  OAI22_X1 U2954 ( .A1(n7258), .A2(n3407), .B1(n3278), .B2(n1376), .ZN(n6128)
         );
  OAI22_X1 U2955 ( .A1(n3129), .A2(n3407), .B1(n3278), .B2(n1375), .ZN(n6129)
         );
  OAI22_X1 U2956 ( .A1(n3119), .A2(n3407), .B1(n3278), .B2(n1374), .ZN(n6130)
         );
  OAI22_X1 U2957 ( .A1(n3116), .A2(n3407), .B1(n3278), .B2(n1373), .ZN(n6131)
         );
  OAI22_X1 U2958 ( .A1(n3106), .A2(n3407), .B1(n3278), .B2(n1372), .ZN(n6132)
         );
  OAI22_X1 U2959 ( .A1(n3093), .A2(n3407), .B1(n3278), .B2(n1371), .ZN(n6133)
         );
  OAI22_X1 U2960 ( .A1(n7252), .A2(n3407), .B1(n3278), .B2(n1370), .ZN(n6134)
         );
  OAI22_X1 U2961 ( .A1(n7251), .A2(n3407), .B1(n3278), .B2(n1369), .ZN(n6135)
         );
  OAI22_X1 U2962 ( .A1(n7258), .A2(n3408), .B1(n7226), .B2(n1368), .ZN(n6136)
         );
  OAI22_X1 U2963 ( .A1(n3128), .A2(n3408), .B1(n7226), .B2(n1367), .ZN(n6137)
         );
  OAI22_X1 U2964 ( .A1(n3119), .A2(n3408), .B1(n7226), .B2(n1366), .ZN(n6138)
         );
  OAI22_X1 U2965 ( .A1(n7255), .A2(n3408), .B1(n7226), .B2(n1365), .ZN(n6139)
         );
  OAI22_X1 U2966 ( .A1(n3100), .A2(n3408), .B1(n7226), .B2(n1364), .ZN(n6140)
         );
  OAI22_X1 U2967 ( .A1(n3091), .A2(n3408), .B1(n7226), .B2(n1363), .ZN(n6141)
         );
  OAI22_X1 U2968 ( .A1(n7252), .A2(n3408), .B1(n7226), .B2(n1362), .ZN(n6142)
         );
  OAI22_X1 U2969 ( .A1(n7251), .A2(n3408), .B1(n7226), .B2(n1361), .ZN(n6143)
         );
  OAI22_X1 U2970 ( .A1(n3141), .A2(n3409), .B1(n3342), .B2(n1344), .ZN(n6144)
         );
  OAI22_X1 U2971 ( .A1(n3131), .A2(n3409), .B1(n3342), .B2(n1343), .ZN(n6145)
         );
  OAI22_X1 U2972 ( .A1(n3119), .A2(n3409), .B1(n3342), .B2(n1342), .ZN(n6146)
         );
  OAI22_X1 U2973 ( .A1(n3115), .A2(n3409), .B1(n3342), .B2(n1341), .ZN(n6147)
         );
  OAI22_X1 U2974 ( .A1(n3106), .A2(n3409), .B1(n3342), .B2(n1340), .ZN(n6148)
         );
  OAI22_X1 U2975 ( .A1(n3098), .A2(n3409), .B1(n3342), .B2(n1339), .ZN(n6149)
         );
  OAI22_X1 U2976 ( .A1(n3090), .A2(n3409), .B1(n3342), .B2(n1338), .ZN(n6150)
         );
  OAI22_X1 U2977 ( .A1(n3081), .A2(n3409), .B1(n3342), .B2(n1337), .ZN(n6151)
         );
  OAI22_X1 U2978 ( .A1(n3137), .A2(n3410), .B1(n7162), .B2(n1336), .ZN(n6152)
         );
  OAI22_X1 U2979 ( .A1(n3129), .A2(n3410), .B1(n7162), .B2(n1335), .ZN(n6153)
         );
  OAI22_X1 U2980 ( .A1(n3118), .A2(n3410), .B1(n7162), .B2(n1334), .ZN(n6154)
         );
  OAI22_X1 U2981 ( .A1(n3112), .A2(n3410), .B1(n7162), .B2(n1333), .ZN(n6155)
         );
  OAI22_X1 U2982 ( .A1(n3106), .A2(n3410), .B1(n7162), .B2(n1332), .ZN(n6156)
         );
  OAI22_X1 U2983 ( .A1(n3093), .A2(n3410), .B1(n7162), .B2(n1331), .ZN(n6157)
         );
  OAI22_X1 U2984 ( .A1(n3090), .A2(n3410), .B1(n7162), .B2(n1330), .ZN(n6158)
         );
  OAI22_X1 U2985 ( .A1(n3081), .A2(n3410), .B1(n7162), .B2(n1329), .ZN(n6159)
         );
  OAI22_X1 U2986 ( .A1(n3140), .A2(n3411), .B1(n3262), .B2(n1312), .ZN(n6160)
         );
  OAI22_X1 U2987 ( .A1(n3129), .A2(n3411), .B1(n3262), .B2(n1311), .ZN(n6161)
         );
  OAI22_X1 U2988 ( .A1(n3118), .A2(n3411), .B1(n3262), .B2(n1310), .ZN(n6162)
         );
  OAI22_X1 U2989 ( .A1(n3111), .A2(n3411), .B1(n3262), .B2(n1309), .ZN(n6163)
         );
  OAI22_X1 U2990 ( .A1(n7254), .A2(n3411), .B1(n3262), .B2(n1308), .ZN(n6164)
         );
  OAI22_X1 U2991 ( .A1(n3099), .A2(n3411), .B1(n3262), .B2(n1307), .ZN(n6165)
         );
  OAI22_X1 U2992 ( .A1(n3086), .A2(n3411), .B1(n3262), .B2(n1306), .ZN(n6166)
         );
  OAI22_X1 U2993 ( .A1(n3077), .A2(n3411), .B1(n3262), .B2(n1305), .ZN(n6167)
         );
  OAI22_X1 U2994 ( .A1(n3139), .A2(n3412), .B1(n7210), .B2(n1304), .ZN(n6168)
         );
  OAI22_X1 U2995 ( .A1(n3136), .A2(n3412), .B1(n7210), .B2(n1303), .ZN(n6169)
         );
  OAI22_X1 U2996 ( .A1(n3119), .A2(n3412), .B1(n7210), .B2(n1302), .ZN(n6170)
         );
  OAI22_X1 U2997 ( .A1(n3113), .A2(n3412), .B1(n7210), .B2(n1301), .ZN(n6171)
         );
  OAI22_X1 U2998 ( .A1(n3104), .A2(n3412), .B1(n7210), .B2(n1300), .ZN(n6172)
         );
  OAI22_X1 U2999 ( .A1(n3091), .A2(n3412), .B1(n7210), .B2(n1299), .ZN(n6173)
         );
  OAI22_X1 U3000 ( .A1(n3084), .A2(n3412), .B1(n7210), .B2(n1298), .ZN(n6174)
         );
  OAI22_X1 U3001 ( .A1(n3075), .A2(n3412), .B1(n7210), .B2(n1297), .ZN(n6175)
         );
  OAI22_X1 U3002 ( .A1(n3142), .A2(n3413), .B1(n3326), .B2(n1280), .ZN(n6176)
         );
  OAI22_X1 U3003 ( .A1(n3135), .A2(n3413), .B1(n3326), .B2(n1279), .ZN(n6177)
         );
  OAI22_X1 U3004 ( .A1(n3118), .A2(n3413), .B1(n3326), .B2(n1278), .ZN(n6178)
         );
  OAI22_X1 U3005 ( .A1(n3111), .A2(n3413), .B1(n3326), .B2(n1277), .ZN(n6179)
         );
  OAI22_X1 U3006 ( .A1(n3101), .A2(n3413), .B1(n3326), .B2(n1276), .ZN(n6180)
         );
  OAI22_X1 U3007 ( .A1(n3093), .A2(n3413), .B1(n3326), .B2(n1275), .ZN(n6181)
         );
  OAI22_X1 U3008 ( .A1(n3090), .A2(n3413), .B1(n3326), .B2(n1274), .ZN(n6182)
         );
  OAI22_X1 U3009 ( .A1(n3081), .A2(n3413), .B1(n3326), .B2(n1273), .ZN(n6183)
         );
  OAI22_X1 U3010 ( .A1(n3137), .A2(n3414), .B1(n7146), .B2(n1272), .ZN(n6184)
         );
  OAI22_X1 U3011 ( .A1(n3136), .A2(n3414), .B1(n7146), .B2(n1271), .ZN(n6185)
         );
  OAI22_X1 U3012 ( .A1(n3118), .A2(n3414), .B1(n7146), .B2(n1270), .ZN(n6186)
         );
  OAI22_X1 U3013 ( .A1(n3112), .A2(n3414), .B1(n7146), .B2(n1269), .ZN(n6187)
         );
  OAI22_X1 U3014 ( .A1(n3107), .A2(n3414), .B1(n7146), .B2(n1268), .ZN(n6188)
         );
  OAI22_X1 U3015 ( .A1(n3091), .A2(n3414), .B1(n7146), .B2(n1267), .ZN(n6189)
         );
  OAI22_X1 U3016 ( .A1(n3087), .A2(n3414), .B1(n7146), .B2(n1266), .ZN(n6190)
         );
  OAI22_X1 U3017 ( .A1(n3078), .A2(n3414), .B1(n7146), .B2(n1265), .ZN(n6191)
         );
  OAI22_X1 U3018 ( .A1(n3140), .A2(n3415), .B1(n3246), .B2(n1248), .ZN(n6192)
         );
  OAI22_X1 U3019 ( .A1(n3134), .A2(n3415), .B1(n3246), .B2(n1247), .ZN(n6193)
         );
  OAI22_X1 U3020 ( .A1(n3118), .A2(n3415), .B1(n3246), .B2(n1246), .ZN(n6194)
         );
  OAI22_X1 U3021 ( .A1(n3111), .A2(n3415), .B1(n3246), .B2(n1245), .ZN(n6195)
         );
  OAI22_X1 U3022 ( .A1(n3104), .A2(n3415), .B1(n3246), .B2(n1244), .ZN(n6196)
         );
  OAI22_X1 U3023 ( .A1(n3095), .A2(n3415), .B1(n3246), .B2(n1243), .ZN(n6197)
         );
  OAI22_X1 U3024 ( .A1(n3084), .A2(n3415), .B1(n3246), .B2(n1242), .ZN(n6198)
         );
  OAI22_X1 U3025 ( .A1(n3075), .A2(n3415), .B1(n3246), .B2(n1241), .ZN(n6199)
         );
  OAI22_X1 U3026 ( .A1(n3139), .A2(n3416), .B1(n7194), .B2(n1240), .ZN(n6200)
         );
  OAI22_X1 U3027 ( .A1(n3133), .A2(n3416), .B1(n7194), .B2(n1239), .ZN(n6201)
         );
  OAI22_X1 U3028 ( .A1(n3119), .A2(n3416), .B1(n7194), .B2(n1238), .ZN(n6202)
         );
  OAI22_X1 U3029 ( .A1(n3117), .A2(n3416), .B1(n7194), .B2(n1237), .ZN(n6203)
         );
  OAI22_X1 U3030 ( .A1(n3101), .A2(n3416), .B1(n7194), .B2(n1236), .ZN(n6204)
         );
  OAI22_X1 U3031 ( .A1(n7253), .A2(n3416), .B1(n7194), .B2(n1235), .ZN(n6205)
         );
  OAI22_X1 U3032 ( .A1(n3085), .A2(n3416), .B1(n7194), .B2(n1234), .ZN(n6206)
         );
  OAI22_X1 U3033 ( .A1(n3076), .A2(n3416), .B1(n7194), .B2(n1233), .ZN(n6207)
         );
  OAI22_X1 U3034 ( .A1(n3144), .A2(n3419), .B1(n3310), .B2(n1216), .ZN(n6208)
         );
  OAI22_X1 U3035 ( .A1(n3132), .A2(n3419), .B1(n3310), .B2(n1215), .ZN(n6209)
         );
  OAI22_X1 U3036 ( .A1(n3118), .A2(n3419), .B1(n3310), .B2(n1214), .ZN(n6210)
         );
  OAI22_X1 U3037 ( .A1(n3114), .A2(n3419), .B1(n3310), .B2(n1213), .ZN(n6211)
         );
  OAI22_X1 U3038 ( .A1(n3101), .A2(n3419), .B1(n3310), .B2(n1212), .ZN(n6212)
         );
  OAI22_X1 U3039 ( .A1(n3095), .A2(n3419), .B1(n3310), .B2(n1211), .ZN(n6213)
         );
  OAI22_X1 U3040 ( .A1(n3090), .A2(n3419), .B1(n3310), .B2(n1210), .ZN(n6214)
         );
  OAI22_X1 U3041 ( .A1(n3081), .A2(n3419), .B1(n3310), .B2(n1209), .ZN(n6215)
         );
  OAI22_X1 U3042 ( .A1(n3137), .A2(n3421), .B1(n7130), .B2(n1208), .ZN(n6216)
         );
  OAI22_X1 U3043 ( .A1(n3131), .A2(n3421), .B1(n7130), .B2(n1207), .ZN(n6217)
         );
  OAI22_X1 U3044 ( .A1(n3119), .A2(n3421), .B1(n7130), .B2(n1206), .ZN(n6218)
         );
  OAI22_X1 U3045 ( .A1(n3117), .A2(n3421), .B1(n7130), .B2(n1205), .ZN(n6219)
         );
  OAI22_X1 U3046 ( .A1(n3104), .A2(n3421), .B1(n7130), .B2(n1204), .ZN(n6220)
         );
  OAI22_X1 U3047 ( .A1(n3091), .A2(n3421), .B1(n7130), .B2(n1203), .ZN(n6221)
         );
  OAI22_X1 U3048 ( .A1(n7252), .A2(n3421), .B1(n7130), .B2(n1202), .ZN(n6222)
         );
  OAI22_X1 U3049 ( .A1(n7251), .A2(n3421), .B1(n7130), .B2(n1201), .ZN(n6223)
         );
  OAI22_X1 U3050 ( .A1(n3140), .A2(n3422), .B1(n3293), .B2(n1184), .ZN(n6224)
         );
  OAI22_X1 U3051 ( .A1(n3133), .A2(n3422), .B1(n3293), .B2(n1183), .ZN(n6225)
         );
  OAI22_X1 U3052 ( .A1(n3120), .A2(n3422), .B1(n3293), .B2(n1182), .ZN(n6226)
         );
  OAI22_X1 U3053 ( .A1(n3111), .A2(n3422), .B1(n3293), .B2(n1181), .ZN(n6227)
         );
  OAI22_X1 U3054 ( .A1(n3101), .A2(n3422), .B1(n3293), .B2(n1180), .ZN(n6228)
         );
  OAI22_X1 U3055 ( .A1(n3098), .A2(n3422), .B1(n3293), .B2(n1179), .ZN(n6229)
         );
  OAI22_X1 U3056 ( .A1(n3085), .A2(n3422), .B1(n3293), .B2(n1178), .ZN(n6230)
         );
  OAI22_X1 U3057 ( .A1(n3076), .A2(n3422), .B1(n3293), .B2(n1177), .ZN(n6231)
         );
  OAI22_X1 U3058 ( .A1(n3139), .A2(n3423), .B1(n7241), .B2(n1176), .ZN(n6232)
         );
  OAI22_X1 U3059 ( .A1(n3131), .A2(n3423), .B1(n7241), .B2(n1175), .ZN(n6233)
         );
  OAI22_X1 U3060 ( .A1(n3119), .A2(n3423), .B1(n7241), .B2(n1174), .ZN(n6234)
         );
  OAI22_X1 U3061 ( .A1(n3115), .A2(n3423), .B1(n7241), .B2(n1173), .ZN(n6235)
         );
  OAI22_X1 U3062 ( .A1(n3104), .A2(n3423), .B1(n7241), .B2(n1172), .ZN(n6236)
         );
  OAI22_X1 U3063 ( .A1(n3091), .A2(n3423), .B1(n7241), .B2(n1171), .ZN(n6237)
         );
  OAI22_X1 U3064 ( .A1(n3084), .A2(n3423), .B1(n7241), .B2(n1170), .ZN(n6238)
         );
  OAI22_X1 U3065 ( .A1(n3075), .A2(n3423), .B1(n7241), .B2(n1169), .ZN(n6239)
         );
  OAI22_X1 U3066 ( .A1(n3142), .A2(n3424), .B1(n7112), .B2(n1152), .ZN(n6240)
         );
  OAI22_X1 U3067 ( .A1(n3132), .A2(n3424), .B1(n7112), .B2(n1151), .ZN(n6241)
         );
  OAI22_X1 U3068 ( .A1(n3118), .A2(n3424), .B1(n7112), .B2(n1150), .ZN(n6242)
         );
  OAI22_X1 U3069 ( .A1(n7255), .A2(n3424), .B1(n7112), .B2(n1149), .ZN(n6243)
         );
  OAI22_X1 U3070 ( .A1(n3104), .A2(n3424), .B1(n7112), .B2(n1148), .ZN(n6244)
         );
  OAI22_X1 U3071 ( .A1(n3099), .A2(n3424), .B1(n7112), .B2(n1147), .ZN(n6245)
         );
  OAI22_X1 U3072 ( .A1(n3084), .A2(n3424), .B1(n7112), .B2(n1146), .ZN(n6246)
         );
  OAI22_X1 U3073 ( .A1(n3075), .A2(n3424), .B1(n7112), .B2(n1145), .ZN(n6247)
         );
  OAI22_X1 U3074 ( .A1(n3139), .A2(n3425), .B1(n7177), .B2(n1144), .ZN(n6248)
         );
  OAI22_X1 U3075 ( .A1(n7257), .A2(n3425), .B1(n7177), .B2(n1143), .ZN(n6249)
         );
  OAI22_X1 U3076 ( .A1(n3120), .A2(n3425), .B1(n7177), .B2(n1142), .ZN(n6250)
         );
  OAI22_X1 U3077 ( .A1(n3111), .A2(n3425), .B1(n7177), .B2(n1141), .ZN(n6251)
         );
  OAI22_X1 U3078 ( .A1(n3100), .A2(n3425), .B1(n7177), .B2(n1140), .ZN(n6252)
         );
  OAI22_X1 U3079 ( .A1(n3091), .A2(n3425), .B1(n7177), .B2(n1139), .ZN(n6253)
         );
  OAI22_X1 U3080 ( .A1(n3086), .A2(n3425), .B1(n7177), .B2(n1138), .ZN(n6254)
         );
  OAI22_X1 U3081 ( .A1(n3077), .A2(n3425), .B1(n7177), .B2(n1137), .ZN(n6255)
         );
  OAI22_X1 U3082 ( .A1(n3143), .A2(n3426), .B1(n3277), .B2(n1120), .ZN(n6256)
         );
  OAI22_X1 U3083 ( .A1(n3128), .A2(n3426), .B1(n3277), .B2(n1119), .ZN(n6257)
         );
  OAI22_X1 U3084 ( .A1(n3120), .A2(n3426), .B1(n3277), .B2(n1118), .ZN(n6258)
         );
  OAI22_X1 U3085 ( .A1(n3112), .A2(n3426), .B1(n3277), .B2(n1117), .ZN(n6259)
         );
  OAI22_X1 U3086 ( .A1(n3100), .A2(n3426), .B1(n3277), .B2(n1116), .ZN(n6260)
         );
  OAI22_X1 U3087 ( .A1(n3092), .A2(n3426), .B1(n3277), .B2(n1115), .ZN(n6261)
         );
  OAI22_X1 U3088 ( .A1(n3084), .A2(n3426), .B1(n3277), .B2(n1114), .ZN(n6262)
         );
  OAI22_X1 U3089 ( .A1(n3075), .A2(n3426), .B1(n3277), .B2(n1113), .ZN(n6263)
         );
  OAI22_X1 U3090 ( .A1(n3137), .A2(n3427), .B1(n7225), .B2(n1112), .ZN(n6264)
         );
  OAI22_X1 U3091 ( .A1(n3134), .A2(n3427), .B1(n7225), .B2(n1111), .ZN(n6265)
         );
  OAI22_X1 U3092 ( .A1(n3120), .A2(n3427), .B1(n7225), .B2(n1110), .ZN(n6266)
         );
  OAI22_X1 U3093 ( .A1(n3111), .A2(n3427), .B1(n7225), .B2(n1109), .ZN(n6267)
         );
  OAI22_X1 U3094 ( .A1(n3107), .A2(n3427), .B1(n7225), .B2(n1108), .ZN(n6268)
         );
  OAI22_X1 U3095 ( .A1(n3092), .A2(n3427), .B1(n7225), .B2(n1107), .ZN(n6269)
         );
  OAI22_X1 U3096 ( .A1(n3090), .A2(n3427), .B1(n7225), .B2(n1106), .ZN(n6270)
         );
  OAI22_X1 U3097 ( .A1(n3081), .A2(n3427), .B1(n7225), .B2(n1105), .ZN(n6271)
         );
  OAI22_X1 U3098 ( .A1(n3139), .A2(n3428), .B1(n3341), .B2(n1088), .ZN(n6272)
         );
  OAI22_X1 U3099 ( .A1(n3129), .A2(n3428), .B1(n3341), .B2(n1087), .ZN(n6273)
         );
  OAI22_X1 U3100 ( .A1(n3121), .A2(n3428), .B1(n3341), .B2(n1086), .ZN(n6274)
         );
  OAI22_X1 U3101 ( .A1(n3113), .A2(n3428), .B1(n3341), .B2(n1085), .ZN(n6275)
         );
  OAI22_X1 U3102 ( .A1(n3100), .A2(n3428), .B1(n3341), .B2(n1084), .ZN(n6276)
         );
  OAI22_X1 U3103 ( .A1(n3092), .A2(n3428), .B1(n3341), .B2(n1083), .ZN(n6277)
         );
  OAI22_X1 U3104 ( .A1(n3087), .A2(n3428), .B1(n3341), .B2(n1082), .ZN(n6278)
         );
  OAI22_X1 U3105 ( .A1(n3078), .A2(n3428), .B1(n3341), .B2(n1081), .ZN(n6279)
         );
  OAI22_X1 U3106 ( .A1(n3140), .A2(n3429), .B1(n7161), .B2(n1080), .ZN(n6280)
         );
  OAI22_X1 U3107 ( .A1(n3128), .A2(n3429), .B1(n7161), .B2(n1079), .ZN(n6281)
         );
  OAI22_X1 U3108 ( .A1(n3118), .A2(n3429), .B1(n7161), .B2(n1078), .ZN(n6282)
         );
  OAI22_X1 U3109 ( .A1(n3111), .A2(n3429), .B1(n7161), .B2(n1077), .ZN(n6283)
         );
  OAI22_X1 U3110 ( .A1(n3100), .A2(n3429), .B1(n7161), .B2(n1076), .ZN(n6284)
         );
  OAI22_X1 U3111 ( .A1(n3092), .A2(n3429), .B1(n7161), .B2(n1075), .ZN(n6285)
         );
  OAI22_X1 U3112 ( .A1(n3084), .A2(n3429), .B1(n7161), .B2(n1074), .ZN(n6286)
         );
  OAI22_X1 U3113 ( .A1(n3075), .A2(n3429), .B1(n7161), .B2(n1073), .ZN(n6287)
         );
  OAI22_X1 U3114 ( .A1(n3145), .A2(n3430), .B1(n3261), .B2(n1056), .ZN(n6288)
         );
  OAI22_X1 U3115 ( .A1(n3135), .A2(n3430), .B1(n3261), .B2(n1055), .ZN(n6289)
         );
  OAI22_X1 U3116 ( .A1(n3120), .A2(n3430), .B1(n3261), .B2(n1054), .ZN(n6290)
         );
  OAI22_X1 U3117 ( .A1(n3115), .A2(n3430), .B1(n3261), .B2(n1053), .ZN(n6291)
         );
  OAI22_X1 U3118 ( .A1(n3104), .A2(n3430), .B1(n3261), .B2(n1052), .ZN(n6292)
         );
  OAI22_X1 U3119 ( .A1(n3092), .A2(n3430), .B1(n3261), .B2(n1051), .ZN(n6293)
         );
  OAI22_X1 U3120 ( .A1(n3090), .A2(n3430), .B1(n3261), .B2(n1050), .ZN(n6294)
         );
  OAI22_X1 U3121 ( .A1(n3081), .A2(n3430), .B1(n3261), .B2(n1049), .ZN(n6295)
         );
  OAI22_X1 U3122 ( .A1(n3137), .A2(n3431), .B1(n7209), .B2(n1048), .ZN(n6296)
         );
  OAI22_X1 U3123 ( .A1(n3129), .A2(n3431), .B1(n7209), .B2(n1047), .ZN(n6297)
         );
  OAI22_X1 U3124 ( .A1(n3118), .A2(n3431), .B1(n7209), .B2(n1046), .ZN(n6298)
         );
  OAI22_X1 U3125 ( .A1(n3111), .A2(n3431), .B1(n7209), .B2(n1045), .ZN(n6299)
         );
  OAI22_X1 U3126 ( .A1(n7254), .A2(n3431), .B1(n7209), .B2(n1044), .ZN(n6300)
         );
  OAI22_X1 U3127 ( .A1(n3092), .A2(n3431), .B1(n7209), .B2(n1043), .ZN(n6301)
         );
  OAI22_X1 U3128 ( .A1(n3088), .A2(n3431), .B1(n7209), .B2(n1042), .ZN(n6302)
         );
  OAI22_X1 U3129 ( .A1(n3079), .A2(n3431), .B1(n7209), .B2(n1041), .ZN(n6303)
         );
  OAI22_X1 U3130 ( .A1(n3139), .A2(n3432), .B1(n3325), .B2(n1024), .ZN(n6304)
         );
  OAI22_X1 U3131 ( .A1(n3136), .A2(n3432), .B1(n3325), .B2(n1023), .ZN(n6305)
         );
  OAI22_X1 U3132 ( .A1(n3120), .A2(n3432), .B1(n3325), .B2(n1022), .ZN(n6306)
         );
  OAI22_X1 U3133 ( .A1(n3114), .A2(n3432), .B1(n3325), .B2(n1021), .ZN(n6307)
         );
  OAI22_X1 U3134 ( .A1(n3101), .A2(n3432), .B1(n3325), .B2(n1020), .ZN(n6308)
         );
  OAI22_X1 U3135 ( .A1(n3092), .A2(n3432), .B1(n3325), .B2(n1019), .ZN(n6309)
         );
  OAI22_X1 U3136 ( .A1(n3084), .A2(n3432), .B1(n3325), .B2(n1018), .ZN(n6310)
         );
  OAI22_X1 U3137 ( .A1(n3075), .A2(n3432), .B1(n3325), .B2(n1017), .ZN(n6311)
         );
  OAI22_X1 U3138 ( .A1(n3140), .A2(n3433), .B1(n7145), .B2(n1016), .ZN(n6312)
         );
  OAI22_X1 U3139 ( .A1(n3128), .A2(n3433), .B1(n7145), .B2(n1015), .ZN(n6313)
         );
  OAI22_X1 U3140 ( .A1(n3120), .A2(n3433), .B1(n7145), .B2(n1014), .ZN(n6314)
         );
  OAI22_X1 U3141 ( .A1(n3111), .A2(n3433), .B1(n7145), .B2(n1013), .ZN(n6315)
         );
  OAI22_X1 U3142 ( .A1(n3100), .A2(n3433), .B1(n7145), .B2(n1012), .ZN(n6316)
         );
  OAI22_X1 U3143 ( .A1(n3092), .A2(n3433), .B1(n7145), .B2(n1011), .ZN(n6317)
         );
  OAI22_X1 U3144 ( .A1(n3090), .A2(n3433), .B1(n7145), .B2(n1010), .ZN(n6318)
         );
  OAI22_X1 U3145 ( .A1(n3081), .A2(n3433), .B1(n7145), .B2(n1009), .ZN(n6319)
         );
  OAI22_X1 U3146 ( .A1(n3141), .A2(n3434), .B1(n3245), .B2(n992), .ZN(n6320)
         );
  OAI22_X1 U3147 ( .A1(n3134), .A2(n3434), .B1(n3245), .B2(n991), .ZN(n6321)
         );
  OAI22_X1 U3148 ( .A1(n3118), .A2(n3434), .B1(n3245), .B2(n990), .ZN(n6322)
         );
  OAI22_X1 U3149 ( .A1(n3115), .A2(n3434), .B1(n3245), .B2(n989), .ZN(n6323)
         );
  OAI22_X1 U3150 ( .A1(n3101), .A2(n3434), .B1(n3245), .B2(n988), .ZN(n6324)
         );
  OAI22_X1 U3151 ( .A1(n3092), .A2(n3434), .B1(n3245), .B2(n987), .ZN(n6325)
         );
  OAI22_X1 U3152 ( .A1(n3089), .A2(n3434), .B1(n3245), .B2(n986), .ZN(n6326)
         );
  OAI22_X1 U3153 ( .A1(n3080), .A2(n3434), .B1(n3245), .B2(n985), .ZN(n6327)
         );
  OAI22_X1 U3154 ( .A1(n3137), .A2(n3435), .B1(n7193), .B2(n984), .ZN(n6328)
         );
  OAI22_X1 U3155 ( .A1(n3129), .A2(n3435), .B1(n7193), .B2(n983), .ZN(n6329)
         );
  OAI22_X1 U3156 ( .A1(n3119), .A2(n3435), .B1(n7193), .B2(n982), .ZN(n6330)
         );
  OAI22_X1 U3157 ( .A1(n3111), .A2(n3435), .B1(n7193), .B2(n981), .ZN(n6331)
         );
  OAI22_X1 U3158 ( .A1(n3108), .A2(n3435), .B1(n7193), .B2(n980), .ZN(n6332)
         );
  OAI22_X1 U3159 ( .A1(n3092), .A2(n3435), .B1(n7193), .B2(n979), .ZN(n6333)
         );
  OAI22_X1 U3160 ( .A1(n3084), .A2(n3435), .B1(n7193), .B2(n978), .ZN(n6334)
         );
  OAI22_X1 U3161 ( .A1(n3075), .A2(n3435), .B1(n7193), .B2(n977), .ZN(n6335)
         );
  OAI22_X1 U3162 ( .A1(n3139), .A2(n3437), .B1(n3309), .B2(n960), .ZN(n6336)
         );
  OAI22_X1 U3163 ( .A1(n3133), .A2(n3437), .B1(n3309), .B2(n959), .ZN(n6337)
         );
  OAI22_X1 U3164 ( .A1(n7256), .A2(n3437), .B1(n3309), .B2(n958), .ZN(n6338)
         );
  OAI22_X1 U3165 ( .A1(n3112), .A2(n3437), .B1(n3309), .B2(n957), .ZN(n6339)
         );
  OAI22_X1 U3166 ( .A1(n3100), .A2(n3437), .B1(n3309), .B2(n956), .ZN(n6340)
         );
  OAI22_X1 U3167 ( .A1(n3092), .A2(n3437), .B1(n3309), .B2(n955), .ZN(n6341)
         );
  OAI22_X1 U3168 ( .A1(n3090), .A2(n3437), .B1(n3309), .B2(n954), .ZN(n6342)
         );
  OAI22_X1 U3169 ( .A1(n3081), .A2(n3437), .B1(n3309), .B2(n953), .ZN(n6343)
         );
  OAI22_X1 U3170 ( .A1(n3140), .A2(n3439), .B1(n7129), .B2(n952), .ZN(n6344)
         );
  OAI22_X1 U3171 ( .A1(n3128), .A2(n3439), .B1(n7129), .B2(n951), .ZN(n6345)
         );
  OAI22_X1 U3172 ( .A1(n7256), .A2(n3439), .B1(n7129), .B2(n950), .ZN(n6346)
         );
  OAI22_X1 U3173 ( .A1(n3111), .A2(n3439), .B1(n7129), .B2(n949), .ZN(n6347)
         );
  OAI22_X1 U3174 ( .A1(n3107), .A2(n3439), .B1(n7129), .B2(n948), .ZN(n6348)
         );
  OAI22_X1 U3175 ( .A1(n3092), .A2(n3439), .B1(n7129), .B2(n947), .ZN(n6349)
         );
  OAI22_X1 U3176 ( .A1(n3085), .A2(n3439), .B1(n7129), .B2(n946), .ZN(n6350)
         );
  OAI22_X1 U3177 ( .A1(n3076), .A2(n3439), .B1(n7129), .B2(n945), .ZN(n6351)
         );
  OAI22_X1 U3178 ( .A1(n3140), .A2(n3440), .B1(n3292), .B2(n928), .ZN(n6352)
         );
  OAI22_X1 U3179 ( .A1(n7257), .A2(n3440), .B1(n3292), .B2(n927), .ZN(n6353)
         );
  OAI22_X1 U3180 ( .A1(n3121), .A2(n3440), .B1(n3292), .B2(n926), .ZN(n6354)
         );
  OAI22_X1 U3181 ( .A1(n3110), .A2(n3440), .B1(n3292), .B2(n925), .ZN(n6355)
         );
  OAI22_X1 U3182 ( .A1(n3102), .A2(n3440), .B1(n3292), .B2(n924), .ZN(n6356)
         );
  OAI22_X1 U3183 ( .A1(n3092), .A2(n3440), .B1(n3292), .B2(n923), .ZN(n6357)
         );
  OAI22_X1 U3184 ( .A1(n3090), .A2(n3440), .B1(n3292), .B2(n922), .ZN(n6358)
         );
  OAI22_X1 U3185 ( .A1(n3081), .A2(n3440), .B1(n3292), .B2(n921), .ZN(n6359)
         );
  OAI22_X1 U3186 ( .A1(n3139), .A2(n3441), .B1(n7240), .B2(n920), .ZN(n6360)
         );
  OAI22_X1 U3187 ( .A1(n3129), .A2(n3441), .B1(n7240), .B2(n919), .ZN(n6361)
         );
  OAI22_X1 U3188 ( .A1(n3121), .A2(n3441), .B1(n7240), .B2(n918), .ZN(n6362)
         );
  OAI22_X1 U3189 ( .A1(n3110), .A2(n3441), .B1(n7240), .B2(n917), .ZN(n6363)
         );
  OAI22_X1 U3190 ( .A1(n3104), .A2(n3441), .B1(n7240), .B2(n916), .ZN(n6364)
         );
  OAI22_X1 U3191 ( .A1(n7253), .A2(n3441), .B1(n7240), .B2(n915), .ZN(n6365)
         );
  OAI22_X1 U3192 ( .A1(n3090), .A2(n3441), .B1(n7240), .B2(n914), .ZN(n6366)
         );
  OAI22_X1 U3193 ( .A1(n3081), .A2(n3441), .B1(n7240), .B2(n913), .ZN(n6367)
         );
  OAI22_X1 U3194 ( .A1(n3139), .A2(n3442), .B1(n7111), .B2(n896), .ZN(n6368)
         );
  OAI22_X1 U3195 ( .A1(n3130), .A2(n3442), .B1(n7111), .B2(n895), .ZN(n6369)
         );
  OAI22_X1 U3196 ( .A1(n3121), .A2(n3442), .B1(n7111), .B2(n894), .ZN(n6370)
         );
  OAI22_X1 U3197 ( .A1(n3110), .A2(n3442), .B1(n7111), .B2(n893), .ZN(n6371)
         );
  OAI22_X1 U3198 ( .A1(n3101), .A2(n3442), .B1(n7111), .B2(n892), .ZN(n6372)
         );
  OAI22_X1 U3199 ( .A1(n7253), .A2(n3442), .B1(n7111), .B2(n891), .ZN(n6373)
         );
  OAI22_X1 U3200 ( .A1(n3090), .A2(n3442), .B1(n7111), .B2(n890), .ZN(n6374)
         );
  OAI22_X1 U3201 ( .A1(n3081), .A2(n3442), .B1(n7111), .B2(n889), .ZN(n6375)
         );
  OAI22_X1 U3202 ( .A1(n3139), .A2(n3443), .B1(n7176), .B2(n888), .ZN(n6376)
         );
  OAI22_X1 U3203 ( .A1(n3128), .A2(n3443), .B1(n7176), .B2(n887), .ZN(n6377)
         );
  OAI22_X1 U3204 ( .A1(n3121), .A2(n3443), .B1(n7176), .B2(n886), .ZN(n6378)
         );
  OAI22_X1 U3205 ( .A1(n3110), .A2(n3443), .B1(n7176), .B2(n885), .ZN(n6379)
         );
  OAI22_X1 U3206 ( .A1(n3108), .A2(n3443), .B1(n7176), .B2(n884), .ZN(n6380)
         );
  OAI22_X1 U3207 ( .A1(n7253), .A2(n3443), .B1(n7176), .B2(n883), .ZN(n6381)
         );
  OAI22_X1 U3208 ( .A1(n3083), .A2(n3443), .B1(n7176), .B2(n882), .ZN(n6382)
         );
  OAI22_X1 U3209 ( .A1(n3074), .A2(n3443), .B1(n7176), .B2(n881), .ZN(n6383)
         );
  OAI22_X1 U3210 ( .A1(n3139), .A2(n3444), .B1(n3276), .B2(n864), .ZN(n6384)
         );
  OAI22_X1 U3211 ( .A1(n3130), .A2(n3444), .B1(n3276), .B2(n863), .ZN(n6385)
         );
  OAI22_X1 U3212 ( .A1(n3121), .A2(n3444), .B1(n3276), .B2(n862), .ZN(n6386)
         );
  OAI22_X1 U3213 ( .A1(n3110), .A2(n3444), .B1(n3276), .B2(n861), .ZN(n6387)
         );
  OAI22_X1 U3214 ( .A1(n3102), .A2(n3444), .B1(n3276), .B2(n860), .ZN(n6388)
         );
  OAI22_X1 U3215 ( .A1(n7253), .A2(n3444), .B1(n3276), .B2(n859), .ZN(n6389)
         );
  OAI22_X1 U3216 ( .A1(n3090), .A2(n3444), .B1(n3276), .B2(n858), .ZN(n6390)
         );
  OAI22_X1 U3217 ( .A1(n3081), .A2(n3444), .B1(n3276), .B2(n857), .ZN(n6391)
         );
  OAI22_X1 U3218 ( .A1(n3139), .A2(n3445), .B1(n7224), .B2(n856), .ZN(n6392)
         );
  OAI22_X1 U3219 ( .A1(n7257), .A2(n3445), .B1(n7224), .B2(n855), .ZN(n6393)
         );
  OAI22_X1 U3220 ( .A1(n3121), .A2(n3445), .B1(n7224), .B2(n854), .ZN(n6394)
         );
  OAI22_X1 U3221 ( .A1(n3110), .A2(n3445), .B1(n7224), .B2(n853), .ZN(n6395)
         );
  OAI22_X1 U3222 ( .A1(n3106), .A2(n3445), .B1(n7224), .B2(n852), .ZN(n6396)
         );
  OAI22_X1 U3223 ( .A1(n7253), .A2(n3445), .B1(n7224), .B2(n851), .ZN(n6397)
         );
  OAI22_X1 U3224 ( .A1(n3082), .A2(n3445), .B1(n7224), .B2(n850), .ZN(n6398)
         );
  OAI22_X1 U3225 ( .A1(n3073), .A2(n3445), .B1(n7224), .B2(n849), .ZN(n6399)
         );
  OAI22_X1 U3226 ( .A1(n3139), .A2(n3446), .B1(n3340), .B2(n832), .ZN(n6400)
         );
  OAI22_X1 U3227 ( .A1(n7257), .A2(n3446), .B1(n3340), .B2(n831), .ZN(n6401)
         );
  OAI22_X1 U3228 ( .A1(n3121), .A2(n3446), .B1(n3340), .B2(n830), .ZN(n6402)
         );
  OAI22_X1 U3229 ( .A1(n3110), .A2(n3446), .B1(n3340), .B2(n829), .ZN(n6403)
         );
  OAI22_X1 U3230 ( .A1(n3107), .A2(n3446), .B1(n3340), .B2(n828), .ZN(n6404)
         );
  OAI22_X1 U3231 ( .A1(n7253), .A2(n3446), .B1(n3340), .B2(n827), .ZN(n6405)
         );
  OAI22_X1 U3232 ( .A1(n3082), .A2(n3446), .B1(n3340), .B2(n826), .ZN(n6406)
         );
  OAI22_X1 U3233 ( .A1(n3073), .A2(n3446), .B1(n3340), .B2(n825), .ZN(n6407)
         );
  OAI22_X1 U3234 ( .A1(n3139), .A2(n3447), .B1(n7160), .B2(n824), .ZN(n6408)
         );
  OAI22_X1 U3235 ( .A1(n7257), .A2(n3447), .B1(n7160), .B2(n823), .ZN(n6409)
         );
  OAI22_X1 U3236 ( .A1(n3121), .A2(n3447), .B1(n7160), .B2(n822), .ZN(n6410)
         );
  OAI22_X1 U3237 ( .A1(n3110), .A2(n3447), .B1(n7160), .B2(n821), .ZN(n6411)
         );
  OAI22_X1 U3238 ( .A1(n3108), .A2(n3447), .B1(n7160), .B2(n820), .ZN(n6412)
         );
  OAI22_X1 U3239 ( .A1(n7253), .A2(n3447), .B1(n7160), .B2(n819), .ZN(n6413)
         );
  OAI22_X1 U3240 ( .A1(n7252), .A2(n3447), .B1(n7160), .B2(n818), .ZN(n6414)
         );
  OAI22_X1 U3241 ( .A1(n7251), .A2(n3447), .B1(n7160), .B2(n817), .ZN(n6415)
         );
  OAI22_X1 U3242 ( .A1(n3139), .A2(n3448), .B1(n3260), .B2(n800), .ZN(n6416)
         );
  OAI22_X1 U3243 ( .A1(n7257), .A2(n3448), .B1(n3260), .B2(n799), .ZN(n6417)
         );
  OAI22_X1 U3244 ( .A1(n3121), .A2(n3448), .B1(n3260), .B2(n798), .ZN(n6418)
         );
  OAI22_X1 U3245 ( .A1(n3110), .A2(n3448), .B1(n3260), .B2(n797), .ZN(n6419)
         );
  OAI22_X1 U3246 ( .A1(n3105), .A2(n3448), .B1(n3260), .B2(n796), .ZN(n6420)
         );
  OAI22_X1 U3247 ( .A1(n7253), .A2(n3448), .B1(n3260), .B2(n795), .ZN(n6421)
         );
  OAI22_X1 U3248 ( .A1(n3083), .A2(n3448), .B1(n3260), .B2(n794), .ZN(n6422)
         );
  OAI22_X1 U3249 ( .A1(n3074), .A2(n3448), .B1(n3260), .B2(n793), .ZN(n6423)
         );
  OAI22_X1 U3250 ( .A1(n3139), .A2(n3449), .B1(n7208), .B2(n792), .ZN(n6424)
         );
  OAI22_X1 U3251 ( .A1(n7257), .A2(n3449), .B1(n7208), .B2(n791), .ZN(n6425)
         );
  OAI22_X1 U3252 ( .A1(n3121), .A2(n3449), .B1(n7208), .B2(n790), .ZN(n6426)
         );
  OAI22_X1 U3253 ( .A1(n3110), .A2(n3449), .B1(n7208), .B2(n789), .ZN(n6427)
         );
  OAI22_X1 U3254 ( .A1(n3104), .A2(n3449), .B1(n7208), .B2(n788), .ZN(n6428)
         );
  OAI22_X1 U3255 ( .A1(n3092), .A2(n3449), .B1(n7208), .B2(n787), .ZN(n6429)
         );
  OAI22_X1 U3256 ( .A1(n7252), .A2(n3449), .B1(n7208), .B2(n786), .ZN(n6430)
         );
  OAI22_X1 U3257 ( .A1(n7251), .A2(n3449), .B1(n7208), .B2(n785), .ZN(n6431)
         );
  OAI22_X1 U3258 ( .A1(n3139), .A2(n3450), .B1(n3324), .B2(n768), .ZN(n6432)
         );
  OAI22_X1 U3259 ( .A1(n7257), .A2(n3450), .B1(n3324), .B2(n767), .ZN(n6433)
         );
  OAI22_X1 U3260 ( .A1(n3121), .A2(n3450), .B1(n3324), .B2(n766), .ZN(n6434)
         );
  OAI22_X1 U3261 ( .A1(n3110), .A2(n3450), .B1(n3324), .B2(n765), .ZN(n6435)
         );
  OAI22_X1 U3262 ( .A1(n3101), .A2(n3450), .B1(n3324), .B2(n764), .ZN(n6436)
         );
  OAI22_X1 U3263 ( .A1(n3092), .A2(n3450), .B1(n3324), .B2(n763), .ZN(n6437)
         );
  OAI22_X1 U3264 ( .A1(n7252), .A2(n3450), .B1(n3324), .B2(n762), .ZN(n6438)
         );
  OAI22_X1 U3265 ( .A1(n7251), .A2(n3450), .B1(n3324), .B2(n761), .ZN(n6439)
         );
  OAI22_X1 U3266 ( .A1(n3139), .A2(n3451), .B1(n7144), .B2(n760), .ZN(n6440)
         );
  OAI22_X1 U3267 ( .A1(n7257), .A2(n3451), .B1(n7144), .B2(n759), .ZN(n6441)
         );
  OAI22_X1 U3268 ( .A1(n3121), .A2(n3451), .B1(n7144), .B2(n758), .ZN(n6442)
         );
  OAI22_X1 U3269 ( .A1(n3110), .A2(n3451), .B1(n7144), .B2(n757), .ZN(n6443)
         );
  OAI22_X1 U3270 ( .A1(n3107), .A2(n3451), .B1(n7144), .B2(n756), .ZN(n6444)
         );
  OAI22_X1 U3271 ( .A1(n3092), .A2(n3451), .B1(n7144), .B2(n755), .ZN(n6445)
         );
  OAI22_X1 U3272 ( .A1(n3086), .A2(n3451), .B1(n7144), .B2(n754), .ZN(n6446)
         );
  OAI22_X1 U3273 ( .A1(n3077), .A2(n3451), .B1(n7144), .B2(n753), .ZN(n6447)
         );
  OAI22_X1 U3274 ( .A1(n3142), .A2(n3452), .B1(n3244), .B2(n736), .ZN(n6448)
         );
  OAI22_X1 U3275 ( .A1(n3128), .A2(n3452), .B1(n3244), .B2(n735), .ZN(n6449)
         );
  OAI22_X1 U3276 ( .A1(n7256), .A2(n3452), .B1(n3244), .B2(n734), .ZN(n6450)
         );
  OAI22_X1 U3277 ( .A1(n3110), .A2(n3452), .B1(n3244), .B2(n733), .ZN(n6451)
         );
  OAI22_X1 U3278 ( .A1(n3102), .A2(n3452), .B1(n3244), .B2(n732), .ZN(n6452)
         );
  OAI22_X1 U3279 ( .A1(n3092), .A2(n3452), .B1(n3244), .B2(n731), .ZN(n6453)
         );
  OAI22_X1 U3280 ( .A1(n3084), .A2(n3452), .B1(n3244), .B2(n730), .ZN(n6454)
         );
  OAI22_X1 U3281 ( .A1(n3075), .A2(n3452), .B1(n3244), .B2(n729), .ZN(n6455)
         );
  OAI22_X1 U3282 ( .A1(n3144), .A2(n3453), .B1(n7192), .B2(n728), .ZN(n6456)
         );
  OAI22_X1 U3283 ( .A1(n3129), .A2(n3453), .B1(n7192), .B2(n727), .ZN(n6457)
         );
  OAI22_X1 U3284 ( .A1(n3127), .A2(n3453), .B1(n7192), .B2(n726), .ZN(n6458)
         );
  OAI22_X1 U3285 ( .A1(n3116), .A2(n3453), .B1(n7192), .B2(n725), .ZN(n6459)
         );
  OAI22_X1 U3286 ( .A1(n3105), .A2(n3453), .B1(n7192), .B2(n724), .ZN(n6460)
         );
  OAI22_X1 U3287 ( .A1(n3099), .A2(n3453), .B1(n7192), .B2(n723), .ZN(n6461)
         );
  OAI22_X1 U3288 ( .A1(n3087), .A2(n3453), .B1(n7192), .B2(n722), .ZN(n6462)
         );
  OAI22_X1 U3289 ( .A1(n3078), .A2(n3453), .B1(n7192), .B2(n721), .ZN(n6463)
         );
  OAI22_X1 U3290 ( .A1(n3143), .A2(n3455), .B1(n3308), .B2(n704), .ZN(n6464)
         );
  OAI22_X1 U3291 ( .A1(n3130), .A2(n3455), .B1(n3308), .B2(n703), .ZN(n6465)
         );
  OAI22_X1 U3292 ( .A1(n3127), .A2(n3455), .B1(n3308), .B2(n702), .ZN(n6466)
         );
  OAI22_X1 U3293 ( .A1(n3109), .A2(n3455), .B1(n3308), .B2(n701), .ZN(n6467)
         );
  OAI22_X1 U3294 ( .A1(n3102), .A2(n3455), .B1(n3308), .B2(n700), .ZN(n6468)
         );
  OAI22_X1 U3295 ( .A1(n3092), .A2(n3455), .B1(n3308), .B2(n699), .ZN(n6469)
         );
  OAI22_X1 U3296 ( .A1(n3088), .A2(n3455), .B1(n3308), .B2(n698), .ZN(n6470)
         );
  OAI22_X1 U3297 ( .A1(n3079), .A2(n3455), .B1(n3308), .B2(n697), .ZN(n6471)
         );
  OAI22_X1 U3298 ( .A1(n3145), .A2(n3457), .B1(n7128), .B2(n696), .ZN(n6472)
         );
  OAI22_X1 U3299 ( .A1(n3129), .A2(n3457), .B1(n7128), .B2(n695), .ZN(n6473)
         );
  OAI22_X1 U3300 ( .A1(n7256), .A2(n3457), .B1(n7128), .B2(n694), .ZN(n6474)
         );
  OAI22_X1 U3301 ( .A1(n3109), .A2(n3457), .B1(n7128), .B2(n693), .ZN(n6475)
         );
  OAI22_X1 U3302 ( .A1(n3103), .A2(n3457), .B1(n7128), .B2(n692), .ZN(n6476)
         );
  OAI22_X1 U3303 ( .A1(n7253), .A2(n3457), .B1(n7128), .B2(n691), .ZN(n6477)
         );
  OAI22_X1 U3304 ( .A1(n3089), .A2(n3457), .B1(n7128), .B2(n690), .ZN(n6478)
         );
  OAI22_X1 U3305 ( .A1(n3080), .A2(n3457), .B1(n7128), .B2(n689), .ZN(n6479)
         );
  OAI22_X1 U3306 ( .A1(n3141), .A2(n3458), .B1(n3291), .B2(n672), .ZN(n6480)
         );
  OAI22_X1 U3307 ( .A1(n3130), .A2(n3458), .B1(n3291), .B2(n671), .ZN(n6481)
         );
  OAI22_X1 U3308 ( .A1(n3118), .A2(n3458), .B1(n3291), .B2(n670), .ZN(n6482)
         );
  OAI22_X1 U3309 ( .A1(n3109), .A2(n3458), .B1(n3291), .B2(n669), .ZN(n6483)
         );
  OAI22_X1 U3310 ( .A1(n3104), .A2(n3458), .B1(n3291), .B2(n668), .ZN(n6484)
         );
  OAI22_X1 U3311 ( .A1(n7253), .A2(n3458), .B1(n3291), .B2(n667), .ZN(n6485)
         );
  OAI22_X1 U3312 ( .A1(n3085), .A2(n3458), .B1(n3291), .B2(n666), .ZN(n6486)
         );
  OAI22_X1 U3313 ( .A1(n3076), .A2(n3458), .B1(n3291), .B2(n665), .ZN(n6487)
         );
  OAI22_X1 U3314 ( .A1(n3142), .A2(n3459), .B1(n7239), .B2(n664), .ZN(n6488)
         );
  OAI22_X1 U3315 ( .A1(n3129), .A2(n3459), .B1(n7239), .B2(n663), .ZN(n6489)
         );
  OAI22_X1 U3316 ( .A1(n3127), .A2(n3459), .B1(n7239), .B2(n662), .ZN(n6490)
         );
  OAI22_X1 U3317 ( .A1(n3109), .A2(n3459), .B1(n7239), .B2(n661), .ZN(n6491)
         );
  OAI22_X1 U3318 ( .A1(n3101), .A2(n3459), .B1(n7239), .B2(n660), .ZN(n6492)
         );
  OAI22_X1 U3319 ( .A1(n7253), .A2(n3459), .B1(n7239), .B2(n659), .ZN(n6493)
         );
  OAI22_X1 U3320 ( .A1(n3086), .A2(n3459), .B1(n7239), .B2(n658), .ZN(n6494)
         );
  OAI22_X1 U3321 ( .A1(n3077), .A2(n3459), .B1(n7239), .B2(n657), .ZN(n6495)
         );
  OAI22_X1 U3322 ( .A1(n3144), .A2(n3460), .B1(n7110), .B2(n640), .ZN(n6496)
         );
  OAI22_X1 U3323 ( .A1(n3130), .A2(n3460), .B1(n7110), .B2(n639), .ZN(n6497)
         );
  OAI22_X1 U3324 ( .A1(n7256), .A2(n3460), .B1(n7110), .B2(n638), .ZN(n6498)
         );
  OAI22_X1 U3325 ( .A1(n3109), .A2(n3460), .B1(n7110), .B2(n637), .ZN(n6499)
         );
  OAI22_X1 U3326 ( .A1(n3108), .A2(n3460), .B1(n7110), .B2(n636), .ZN(n6500)
         );
  OAI22_X1 U3327 ( .A1(n7253), .A2(n3460), .B1(n7110), .B2(n635), .ZN(n6501)
         );
  OAI22_X1 U3328 ( .A1(n3087), .A2(n3460), .B1(n7110), .B2(n634), .ZN(n6502)
         );
  OAI22_X1 U3329 ( .A1(n3078), .A2(n3460), .B1(n7110), .B2(n633), .ZN(n6503)
         );
  OAI22_X1 U3330 ( .A1(n3143), .A2(n3461), .B1(n7175), .B2(n632), .ZN(n6504)
         );
  OAI22_X1 U3331 ( .A1(n3128), .A2(n3461), .B1(n7175), .B2(n631), .ZN(n6505)
         );
  OAI22_X1 U3332 ( .A1(n7256), .A2(n3461), .B1(n7175), .B2(n630), .ZN(n6506)
         );
  OAI22_X1 U3333 ( .A1(n3109), .A2(n3461), .B1(n7175), .B2(n629), .ZN(n6507)
         );
  OAI22_X1 U3334 ( .A1(n3102), .A2(n3461), .B1(n7175), .B2(n628), .ZN(n6508)
         );
  OAI22_X1 U3335 ( .A1(n7253), .A2(n3461), .B1(n7175), .B2(n627), .ZN(n6509)
         );
  OAI22_X1 U3336 ( .A1(n3088), .A2(n3461), .B1(n7175), .B2(n626), .ZN(n6510)
         );
  OAI22_X1 U3337 ( .A1(n3079), .A2(n3461), .B1(n7175), .B2(n625), .ZN(n6511)
         );
  OAI22_X1 U3338 ( .A1(n3145), .A2(n3462), .B1(n3275), .B2(n608), .ZN(n6512)
         );
  OAI22_X1 U3339 ( .A1(n3130), .A2(n3462), .B1(n3275), .B2(n607), .ZN(n6513)
         );
  OAI22_X1 U3340 ( .A1(n3127), .A2(n3462), .B1(n3275), .B2(n606), .ZN(n6514)
         );
  OAI22_X1 U3341 ( .A1(n3109), .A2(n3462), .B1(n3275), .B2(n605), .ZN(n6515)
         );
  OAI22_X1 U3342 ( .A1(n3103), .A2(n3462), .B1(n3275), .B2(n604), .ZN(n6516)
         );
  OAI22_X1 U3343 ( .A1(n7253), .A2(n3462), .B1(n3275), .B2(n603), .ZN(n6517)
         );
  OAI22_X1 U3344 ( .A1(n3089), .A2(n3462), .B1(n3275), .B2(n602), .ZN(n6518)
         );
  OAI22_X1 U3345 ( .A1(n3080), .A2(n3462), .B1(n3275), .B2(n601), .ZN(n6519)
         );
  OAI22_X1 U3346 ( .A1(n3141), .A2(n3463), .B1(n7223), .B2(n600), .ZN(n6520)
         );
  OAI22_X1 U3347 ( .A1(n3129), .A2(n3463), .B1(n7223), .B2(n599), .ZN(n6521)
         );
  OAI22_X1 U3348 ( .A1(n3118), .A2(n3463), .B1(n7223), .B2(n598), .ZN(n6522)
         );
  OAI22_X1 U3349 ( .A1(n3109), .A2(n3463), .B1(n7223), .B2(n597), .ZN(n6523)
         );
  OAI22_X1 U3350 ( .A1(n3105), .A2(n3463), .B1(n7223), .B2(n596), .ZN(n6524)
         );
  OAI22_X1 U3351 ( .A1(n7253), .A2(n3463), .B1(n7223), .B2(n595), .ZN(n6525)
         );
  OAI22_X1 U3352 ( .A1(n3085), .A2(n3463), .B1(n7223), .B2(n594), .ZN(n6526)
         );
  OAI22_X1 U3353 ( .A1(n3076), .A2(n3463), .B1(n7223), .B2(n593), .ZN(n6527)
         );
  OAI22_X1 U3354 ( .A1(n3144), .A2(n3464), .B1(n3339), .B2(n576), .ZN(n6528)
         );
  OAI22_X1 U3355 ( .A1(n3130), .A2(n3464), .B1(n3339), .B2(n575), .ZN(n6529)
         );
  OAI22_X1 U3356 ( .A1(n3122), .A2(n3464), .B1(n3339), .B2(n574), .ZN(n6530)
         );
  OAI22_X1 U3357 ( .A1(n3109), .A2(n3464), .B1(n3339), .B2(n573), .ZN(n6531)
         );
  OAI22_X1 U3358 ( .A1(n3106), .A2(n3464), .B1(n3339), .B2(n572), .ZN(n6532)
         );
  OAI22_X1 U3359 ( .A1(n7253), .A2(n3464), .B1(n3339), .B2(n571), .ZN(n6533)
         );
  OAI22_X1 U3360 ( .A1(n3086), .A2(n3464), .B1(n3339), .B2(n570), .ZN(n6534)
         );
  OAI22_X1 U3361 ( .A1(n3077), .A2(n3464), .B1(n3339), .B2(n569), .ZN(n6535)
         );
  OAI22_X1 U3362 ( .A1(n3143), .A2(n3465), .B1(n7159), .B2(n568), .ZN(n6536)
         );
  OAI22_X1 U3363 ( .A1(n3128), .A2(n3465), .B1(n7159), .B2(n567), .ZN(n6537)
         );
  OAI22_X1 U3364 ( .A1(n7256), .A2(n3465), .B1(n7159), .B2(n566), .ZN(n6538)
         );
  OAI22_X1 U3365 ( .A1(n3114), .A2(n3465), .B1(n7159), .B2(n565), .ZN(n6539)
         );
  OAI22_X1 U3366 ( .A1(n3107), .A2(n3465), .B1(n7159), .B2(n564), .ZN(n6540)
         );
  OAI22_X1 U3367 ( .A1(n7253), .A2(n3465), .B1(n7159), .B2(n563), .ZN(n6541)
         );
  OAI22_X1 U3368 ( .A1(n3087), .A2(n3465), .B1(n7159), .B2(n562), .ZN(n6542)
         );
  OAI22_X1 U3369 ( .A1(n3078), .A2(n3465), .B1(n7159), .B2(n561), .ZN(n6543)
         );
  OAI22_X1 U3370 ( .A1(n3142), .A2(n3466), .B1(n3259), .B2(n560), .ZN(n6544)
         );
  OAI22_X1 U3371 ( .A1(n3130), .A2(n3466), .B1(n3259), .B2(n559), .ZN(n6545)
         );
  OAI22_X1 U3372 ( .A1(n7256), .A2(n3466), .B1(n3259), .B2(n558), .ZN(n6546)
         );
  OAI22_X1 U3373 ( .A1(n3109), .A2(n3466), .B1(n3259), .B2(n557), .ZN(n6547)
         );
  OAI22_X1 U3374 ( .A1(n3108), .A2(n3466), .B1(n3259), .B2(n556), .ZN(n6548)
         );
  OAI22_X1 U3375 ( .A1(n7253), .A2(n3466), .B1(n3259), .B2(n555), .ZN(n6549)
         );
  OAI22_X1 U3376 ( .A1(n3088), .A2(n3466), .B1(n3259), .B2(n554), .ZN(n6550)
         );
  OAI22_X1 U3377 ( .A1(n3079), .A2(n3466), .B1(n3259), .B2(n553), .ZN(n6551)
         );
  OAI22_X1 U3378 ( .A1(n3142), .A2(n3467), .B1(n7207), .B2(n552), .ZN(n6552)
         );
  OAI22_X1 U3379 ( .A1(n3128), .A2(n3467), .B1(n7207), .B2(n551), .ZN(n6553)
         );
  OAI22_X1 U3380 ( .A1(n3120), .A2(n3467), .B1(n7207), .B2(n550), .ZN(n6554)
         );
  OAI22_X1 U3381 ( .A1(n3115), .A2(n3467), .B1(n7207), .B2(n549), .ZN(n6555)
         );
  OAI22_X1 U3382 ( .A1(n3105), .A2(n3467), .B1(n7207), .B2(n548), .ZN(n6556)
         );
  OAI22_X1 U3383 ( .A1(n7253), .A2(n3467), .B1(n7207), .B2(n547), .ZN(n6557)
         );
  OAI22_X1 U3384 ( .A1(n3089), .A2(n3467), .B1(n7207), .B2(n546), .ZN(n6558)
         );
  OAI22_X1 U3385 ( .A1(n3080), .A2(n3467), .B1(n7207), .B2(n545), .ZN(n6559)
         );
  OAI22_X1 U3386 ( .A1(n3141), .A2(n3468), .B1(n3323), .B2(n544), .ZN(n6560)
         );
  OAI22_X1 U3387 ( .A1(n3135), .A2(n3468), .B1(n3323), .B2(n543), .ZN(n6561)
         );
  OAI22_X1 U3388 ( .A1(n3120), .A2(n3468), .B1(n3323), .B2(n542), .ZN(n6562)
         );
  OAI22_X1 U3389 ( .A1(n3110), .A2(n3468), .B1(n3323), .B2(n541), .ZN(n6563)
         );
  OAI22_X1 U3390 ( .A1(n3103), .A2(n3468), .B1(n3323), .B2(n540), .ZN(n6564)
         );
  OAI22_X1 U3391 ( .A1(n3092), .A2(n3468), .B1(n3323), .B2(n539), .ZN(n6565)
         );
  OAI22_X1 U3392 ( .A1(n3086), .A2(n3468), .B1(n3323), .B2(n538), .ZN(n6566)
         );
  OAI22_X1 U3393 ( .A1(n3077), .A2(n3468), .B1(n3323), .B2(n537), .ZN(n6567)
         );
  OAI22_X1 U3394 ( .A1(n7258), .A2(n3469), .B1(n7143), .B2(n536), .ZN(n6568)
         );
  OAI22_X1 U3395 ( .A1(n3129), .A2(n3469), .B1(n7143), .B2(n535), .ZN(n6569)
         );
  OAI22_X1 U3396 ( .A1(n3120), .A2(n3469), .B1(n7143), .B2(n534), .ZN(n6570)
         );
  OAI22_X1 U3397 ( .A1(n3110), .A2(n3469), .B1(n7143), .B2(n533), .ZN(n6571)
         );
  OAI22_X1 U3398 ( .A1(n3102), .A2(n3469), .B1(n7143), .B2(n532), .ZN(n6572)
         );
  OAI22_X1 U3399 ( .A1(n3092), .A2(n3469), .B1(n7143), .B2(n531), .ZN(n6573)
         );
  OAI22_X1 U3400 ( .A1(n3087), .A2(n3469), .B1(n7143), .B2(n530), .ZN(n6574)
         );
  OAI22_X1 U3401 ( .A1(n3078), .A2(n3469), .B1(n7143), .B2(n529), .ZN(n6575)
         );
  OAI22_X1 U3402 ( .A1(n3139), .A2(n3470), .B1(n3243), .B2(n528), .ZN(n6576)
         );
  OAI22_X1 U3403 ( .A1(n7257), .A2(n3470), .B1(n3243), .B2(n527), .ZN(n6577)
         );
  OAI22_X1 U3404 ( .A1(n3121), .A2(n3470), .B1(n3243), .B2(n526), .ZN(n6578)
         );
  OAI22_X1 U3405 ( .A1(n3110), .A2(n3470), .B1(n3243), .B2(n525), .ZN(n6579)
         );
  OAI22_X1 U3406 ( .A1(n3100), .A2(n3470), .B1(n3243), .B2(n524), .ZN(n6580)
         );
  OAI22_X1 U3407 ( .A1(n3094), .A2(n3470), .B1(n3243), .B2(n523), .ZN(n6581)
         );
  OAI22_X1 U3408 ( .A1(n3088), .A2(n3470), .B1(n3243), .B2(n522), .ZN(n6582)
         );
  OAI22_X1 U3409 ( .A1(n3079), .A2(n3470), .B1(n3243), .B2(n521), .ZN(n6583)
         );
  OAI22_X1 U3410 ( .A1(n3145), .A2(n3471), .B1(n7191), .B2(n520), .ZN(n6584)
         );
  OAI22_X1 U3411 ( .A1(n3130), .A2(n3471), .B1(n7191), .B2(n519), .ZN(n6585)
         );
  OAI22_X1 U3412 ( .A1(n3120), .A2(n3471), .B1(n7191), .B2(n518), .ZN(n6586)
         );
  OAI22_X1 U3413 ( .A1(n3110), .A2(n3471), .B1(n7191), .B2(n517), .ZN(n6587)
         );
  OAI22_X1 U3414 ( .A1(n3103), .A2(n3471), .B1(n7191), .B2(n516), .ZN(n6588)
         );
  OAI22_X1 U3415 ( .A1(n3091), .A2(n3471), .B1(n7191), .B2(n515), .ZN(n6589)
         );
  OAI22_X1 U3416 ( .A1(n3089), .A2(n3471), .B1(n7191), .B2(n514), .ZN(n6590)
         );
  OAI22_X1 U3417 ( .A1(n3080), .A2(n3471), .B1(n7191), .B2(n513), .ZN(n6591)
         );
  OAI22_X1 U3418 ( .A1(n3142), .A2(n3472), .B1(n3307), .B2(n512), .ZN(n6592)
         );
  OAI22_X1 U3419 ( .A1(n3130), .A2(n3472), .B1(n3307), .B2(n511), .ZN(n6593)
         );
  OAI22_X1 U3420 ( .A1(n3120), .A2(n3472), .B1(n3307), .B2(n510), .ZN(n6594)
         );
  OAI22_X1 U3421 ( .A1(n3110), .A2(n3472), .B1(n3307), .B2(n509), .ZN(n6595)
         );
  OAI22_X1 U3422 ( .A1(n3100), .A2(n3472), .B1(n3307), .B2(n508), .ZN(n6596)
         );
  OAI22_X1 U3423 ( .A1(n3092), .A2(n3472), .B1(n3307), .B2(n507), .ZN(n6597)
         );
  OAI22_X1 U3424 ( .A1(n3085), .A2(n3472), .B1(n3307), .B2(n506), .ZN(n6598)
         );
  OAI22_X1 U3425 ( .A1(n3076), .A2(n3472), .B1(n3307), .B2(n505), .ZN(n6599)
         );
  OAI22_X1 U3426 ( .A1(n3141), .A2(n3474), .B1(n7127), .B2(n504), .ZN(n6600)
         );
  OAI22_X1 U3427 ( .A1(n3130), .A2(n3474), .B1(n7127), .B2(n503), .ZN(n6601)
         );
  OAI22_X1 U3428 ( .A1(n3120), .A2(n3474), .B1(n7127), .B2(n502), .ZN(n6602)
         );
  OAI22_X1 U3429 ( .A1(n3110), .A2(n3474), .B1(n7127), .B2(n501), .ZN(n6603)
         );
  OAI22_X1 U3430 ( .A1(n3102), .A2(n3474), .B1(n7127), .B2(n500), .ZN(n6604)
         );
  OAI22_X1 U3431 ( .A1(n3091), .A2(n3474), .B1(n7127), .B2(n499), .ZN(n6605)
         );
  OAI22_X1 U3432 ( .A1(n3086), .A2(n3474), .B1(n7127), .B2(n498), .ZN(n6606)
         );
  OAI22_X1 U3433 ( .A1(n3077), .A2(n3474), .B1(n7127), .B2(n497), .ZN(n6607)
         );
  OAI22_X1 U3434 ( .A1(n3144), .A2(n3475), .B1(n3290), .B2(n496), .ZN(n6608)
         );
  OAI22_X1 U3435 ( .A1(n3128), .A2(n3475), .B1(n3290), .B2(n495), .ZN(n6609)
         );
  OAI22_X1 U3436 ( .A1(n3120), .A2(n3475), .B1(n3290), .B2(n494), .ZN(n6610)
         );
  OAI22_X1 U3437 ( .A1(n3110), .A2(n3475), .B1(n3290), .B2(n493), .ZN(n6611)
         );
  OAI22_X1 U3438 ( .A1(n3100), .A2(n3475), .B1(n3290), .B2(n492), .ZN(n6612)
         );
  OAI22_X1 U3439 ( .A1(n3097), .A2(n3475), .B1(n3290), .B2(n491), .ZN(n6613)
         );
  OAI22_X1 U3440 ( .A1(n3087), .A2(n3475), .B1(n3290), .B2(n490), .ZN(n6614)
         );
  OAI22_X1 U3441 ( .A1(n3078), .A2(n3475), .B1(n3290), .B2(n489), .ZN(n6615)
         );
  OAI22_X1 U3442 ( .A1(n3143), .A2(n3476), .B1(n7238), .B2(n488), .ZN(n6616)
         );
  OAI22_X1 U3443 ( .A1(n3129), .A2(n3476), .B1(n7238), .B2(n487), .ZN(n6617)
         );
  OAI22_X1 U3444 ( .A1(n3120), .A2(n3476), .B1(n7238), .B2(n486), .ZN(n6618)
         );
  OAI22_X1 U3445 ( .A1(n3110), .A2(n3476), .B1(n7238), .B2(n485), .ZN(n6619)
         );
  OAI22_X1 U3446 ( .A1(n3105), .A2(n3476), .B1(n7238), .B2(n484), .ZN(n6620)
         );
  OAI22_X1 U3447 ( .A1(n3092), .A2(n3476), .B1(n7238), .B2(n483), .ZN(n6621)
         );
  OAI22_X1 U3448 ( .A1(n3088), .A2(n3476), .B1(n7238), .B2(n482), .ZN(n6622)
         );
  OAI22_X1 U3449 ( .A1(n3079), .A2(n3476), .B1(n7238), .B2(n481), .ZN(n6623)
         );
  OAI22_X1 U3450 ( .A1(n3145), .A2(n3477), .B1(n7109), .B2(n480), .ZN(n6624)
         );
  OAI22_X1 U3451 ( .A1(n3130), .A2(n3477), .B1(n7109), .B2(n479), .ZN(n6625)
         );
  OAI22_X1 U3452 ( .A1(n3120), .A2(n3477), .B1(n7109), .B2(n478), .ZN(n6626)
         );
  OAI22_X1 U3453 ( .A1(n3110), .A2(n3477), .B1(n7109), .B2(n477), .ZN(n6627)
         );
  OAI22_X1 U3454 ( .A1(n3103), .A2(n3477), .B1(n7109), .B2(n476), .ZN(n6628)
         );
  OAI22_X1 U3455 ( .A1(n3092), .A2(n3477), .B1(n7109), .B2(n475), .ZN(n6629)
         );
  OAI22_X1 U3456 ( .A1(n3089), .A2(n3477), .B1(n7109), .B2(n474), .ZN(n6630)
         );
  OAI22_X1 U3457 ( .A1(n3080), .A2(n3477), .B1(n7109), .B2(n473), .ZN(n6631)
         );
  OAI22_X1 U3458 ( .A1(n3142), .A2(n3478), .B1(n7174), .B2(n472), .ZN(n6632)
         );
  OAI22_X1 U3459 ( .A1(n3128), .A2(n3478), .B1(n7174), .B2(n471), .ZN(n6633)
         );
  OAI22_X1 U3460 ( .A1(n3120), .A2(n3478), .B1(n7174), .B2(n470), .ZN(n6634)
         );
  OAI22_X1 U3461 ( .A1(n3110), .A2(n3478), .B1(n7174), .B2(n469), .ZN(n6635)
         );
  OAI22_X1 U3462 ( .A1(n3105), .A2(n3478), .B1(n7174), .B2(n468), .ZN(n6636)
         );
  OAI22_X1 U3463 ( .A1(n7253), .A2(n3478), .B1(n7174), .B2(n467), .ZN(n6637)
         );
  OAI22_X1 U3464 ( .A1(n3085), .A2(n3478), .B1(n7174), .B2(n466), .ZN(n6638)
         );
  OAI22_X1 U3465 ( .A1(n3076), .A2(n3478), .B1(n7174), .B2(n465), .ZN(n6639)
         );
  OAI22_X1 U3466 ( .A1(n3141), .A2(n3479), .B1(n3274), .B2(n464), .ZN(n6640)
         );
  OAI22_X1 U3467 ( .A1(n3130), .A2(n3479), .B1(n3274), .B2(n463), .ZN(n6641)
         );
  OAI22_X1 U3468 ( .A1(n3120), .A2(n3479), .B1(n3274), .B2(n462), .ZN(n6642)
         );
  OAI22_X1 U3469 ( .A1(n3110), .A2(n3479), .B1(n3274), .B2(n461), .ZN(n6643)
         );
  OAI22_X1 U3470 ( .A1(n3106), .A2(n3479), .B1(n3274), .B2(n460), .ZN(n6644)
         );
  OAI22_X1 U3471 ( .A1(n7253), .A2(n3479), .B1(n3274), .B2(n459), .ZN(n6645)
         );
  OAI22_X1 U3472 ( .A1(n3086), .A2(n3479), .B1(n3274), .B2(n458), .ZN(n6646)
         );
  OAI22_X1 U3473 ( .A1(n3077), .A2(n3479), .B1(n3274), .B2(n457), .ZN(n6647)
         );
  OAI22_X1 U3474 ( .A1(n3144), .A2(n3480), .B1(n7222), .B2(n456), .ZN(n6648)
         );
  OAI22_X1 U3475 ( .A1(n3129), .A2(n3480), .B1(n7222), .B2(n455), .ZN(n6649)
         );
  OAI22_X1 U3476 ( .A1(n3120), .A2(n3480), .B1(n7222), .B2(n454), .ZN(n6650)
         );
  OAI22_X1 U3477 ( .A1(n3109), .A2(n3480), .B1(n7222), .B2(n453), .ZN(n6651)
         );
  OAI22_X1 U3478 ( .A1(n3107), .A2(n3480), .B1(n7222), .B2(n452), .ZN(n6652)
         );
  OAI22_X1 U3479 ( .A1(n7253), .A2(n3480), .B1(n7222), .B2(n451), .ZN(n6653)
         );
  OAI22_X1 U3480 ( .A1(n3087), .A2(n3480), .B1(n7222), .B2(n450), .ZN(n6654)
         );
  OAI22_X1 U3481 ( .A1(n3078), .A2(n3480), .B1(n7222), .B2(n449), .ZN(n6655)
         );
  OAI22_X1 U3482 ( .A1(n3137), .A2(n3481), .B1(n3338), .B2(n448), .ZN(n6656)
         );
  OAI22_X1 U3483 ( .A1(n3129), .A2(n3481), .B1(n3338), .B2(n447), .ZN(n6657)
         );
  OAI22_X1 U3484 ( .A1(n7256), .A2(n3481), .B1(n3338), .B2(n446), .ZN(n6658)
         );
  OAI22_X1 U3485 ( .A1(n3117), .A2(n3481), .B1(n3338), .B2(n445), .ZN(n6659)
         );
  OAI22_X1 U3486 ( .A1(n3108), .A2(n3481), .B1(n3338), .B2(n444), .ZN(n6660)
         );
  OAI22_X1 U3487 ( .A1(n7253), .A2(n3481), .B1(n3338), .B2(n443), .ZN(n6661)
         );
  OAI22_X1 U3488 ( .A1(n3088), .A2(n3481), .B1(n3338), .B2(n442), .ZN(n6662)
         );
  OAI22_X1 U3489 ( .A1(n3079), .A2(n3481), .B1(n3338), .B2(n441), .ZN(n6663)
         );
  OAI22_X1 U3490 ( .A1(n3137), .A2(n3482), .B1(n7158), .B2(n440), .ZN(n6664)
         );
  OAI22_X1 U3491 ( .A1(n3129), .A2(n3482), .B1(n7158), .B2(n439), .ZN(n6665)
         );
  OAI22_X1 U3492 ( .A1(n3120), .A2(n3482), .B1(n7158), .B2(n438), .ZN(n6666)
         );
  OAI22_X1 U3493 ( .A1(n3111), .A2(n3482), .B1(n7158), .B2(n437), .ZN(n6667)
         );
  OAI22_X1 U3494 ( .A1(n3100), .A2(n3482), .B1(n7158), .B2(n436), .ZN(n6668)
         );
  OAI22_X1 U3495 ( .A1(n3094), .A2(n3482), .B1(n7158), .B2(n435), .ZN(n6669)
         );
  OAI22_X1 U3496 ( .A1(n3084), .A2(n3482), .B1(n7158), .B2(n434), .ZN(n6670)
         );
  OAI22_X1 U3497 ( .A1(n3075), .A2(n3482), .B1(n7158), .B2(n433), .ZN(n6671)
         );
  OAI22_X1 U3498 ( .A1(n3137), .A2(n3483), .B1(n3258), .B2(n432), .ZN(n6672)
         );
  OAI22_X1 U3499 ( .A1(n3135), .A2(n3483), .B1(n3258), .B2(n431), .ZN(n6673)
         );
  OAI22_X1 U3500 ( .A1(n3121), .A2(n3483), .B1(n3258), .B2(n430), .ZN(n6674)
         );
  OAI22_X1 U3501 ( .A1(n3111), .A2(n3483), .B1(n3258), .B2(n429), .ZN(n6675)
         );
  OAI22_X1 U3502 ( .A1(n3103), .A2(n3483), .B1(n3258), .B2(n428), .ZN(n6676)
         );
  OAI22_X1 U3503 ( .A1(n3099), .A2(n3483), .B1(n3258), .B2(n427), .ZN(n6677)
         );
  OAI22_X1 U3504 ( .A1(n3084), .A2(n3483), .B1(n3258), .B2(n426), .ZN(n6678)
         );
  OAI22_X1 U3505 ( .A1(n3075), .A2(n3483), .B1(n3258), .B2(n425), .ZN(n6679)
         );
  OAI22_X1 U3506 ( .A1(n3137), .A2(n3484), .B1(n7206), .B2(n424), .ZN(n6680)
         );
  OAI22_X1 U3507 ( .A1(n3130), .A2(n3484), .B1(n7206), .B2(n423), .ZN(n6681)
         );
  OAI22_X1 U3508 ( .A1(n7256), .A2(n3484), .B1(n7206), .B2(n422), .ZN(n6682)
         );
  OAI22_X1 U3509 ( .A1(n3111), .A2(n3484), .B1(n7206), .B2(n421), .ZN(n6683)
         );
  OAI22_X1 U3510 ( .A1(n3100), .A2(n3484), .B1(n7206), .B2(n420), .ZN(n6684)
         );
  OAI22_X1 U3511 ( .A1(n3092), .A2(n3484), .B1(n7206), .B2(n419), .ZN(n6685)
         );
  OAI22_X1 U3512 ( .A1(n3084), .A2(n3484), .B1(n7206), .B2(n418), .ZN(n6686)
         );
  OAI22_X1 U3513 ( .A1(n3075), .A2(n3484), .B1(n7206), .B2(n417), .ZN(n6687)
         );
  OAI22_X1 U3514 ( .A1(n3137), .A2(n3485), .B1(n3322), .B2(n416), .ZN(n6688)
         );
  OAI22_X1 U3515 ( .A1(n3128), .A2(n3485), .B1(n3322), .B2(n415), .ZN(n6689)
         );
  OAI22_X1 U3516 ( .A1(n3118), .A2(n3485), .B1(n3322), .B2(n414), .ZN(n6690)
         );
  OAI22_X1 U3517 ( .A1(n3111), .A2(n3485), .B1(n3322), .B2(n413), .ZN(n6691)
         );
  OAI22_X1 U3518 ( .A1(n3102), .A2(n3485), .B1(n3322), .B2(n412), .ZN(n6692)
         );
  OAI22_X1 U3519 ( .A1(n3094), .A2(n3485), .B1(n3322), .B2(n411), .ZN(n6693)
         );
  OAI22_X1 U3520 ( .A1(n3084), .A2(n3485), .B1(n3322), .B2(n410), .ZN(n6694)
         );
  OAI22_X1 U3521 ( .A1(n3075), .A2(n3485), .B1(n3322), .B2(n409), .ZN(n6695)
         );
  OAI22_X1 U3522 ( .A1(n3137), .A2(n3486), .B1(n7142), .B2(n408), .ZN(n6696)
         );
  OAI22_X1 U3523 ( .A1(n3130), .A2(n3486), .B1(n7142), .B2(n407), .ZN(n6697)
         );
  OAI22_X1 U3524 ( .A1(n7256), .A2(n3486), .B1(n7142), .B2(n406), .ZN(n6698)
         );
  OAI22_X1 U3525 ( .A1(n3111), .A2(n3486), .B1(n7142), .B2(n405), .ZN(n6699)
         );
  OAI22_X1 U3526 ( .A1(n3100), .A2(n3486), .B1(n7142), .B2(n404), .ZN(n6700)
         );
  OAI22_X1 U3527 ( .A1(n3094), .A2(n3486), .B1(n7142), .B2(n403), .ZN(n6701)
         );
  OAI22_X1 U3528 ( .A1(n3084), .A2(n3486), .B1(n7142), .B2(n402), .ZN(n6702)
         );
  OAI22_X1 U3529 ( .A1(n3075), .A2(n3486), .B1(n7142), .B2(n401), .ZN(n6703)
         );
  OAI22_X1 U3530 ( .A1(n3137), .A2(n3487), .B1(n3242), .B2(n400), .ZN(n6704)
         );
  OAI22_X1 U3531 ( .A1(n3134), .A2(n3487), .B1(n3242), .B2(n399), .ZN(n6705)
         );
  OAI22_X1 U3532 ( .A1(n3125), .A2(n3487), .B1(n3242), .B2(n398), .ZN(n6706)
         );
  OAI22_X1 U3533 ( .A1(n3111), .A2(n3487), .B1(n3242), .B2(n397), .ZN(n6707)
         );
  OAI22_X1 U3534 ( .A1(n3103), .A2(n3487), .B1(n3242), .B2(n396), .ZN(n6708)
         );
  OAI22_X1 U3535 ( .A1(n3098), .A2(n3487), .B1(n3242), .B2(n395), .ZN(n6709)
         );
  OAI22_X1 U3536 ( .A1(n3084), .A2(n3487), .B1(n3242), .B2(n394), .ZN(n6710)
         );
  OAI22_X1 U3537 ( .A1(n3075), .A2(n3487), .B1(n3242), .B2(n393), .ZN(n6711)
         );
  OAI22_X1 U3538 ( .A1(n3137), .A2(n3488), .B1(n7190), .B2(n392), .ZN(n6712)
         );
  OAI22_X1 U3539 ( .A1(n3130), .A2(n3488), .B1(n7190), .B2(n391), .ZN(n6713)
         );
  OAI22_X1 U3540 ( .A1(n7256), .A2(n3488), .B1(n7190), .B2(n390), .ZN(n6714)
         );
  OAI22_X1 U3541 ( .A1(n3111), .A2(n3488), .B1(n7190), .B2(n389), .ZN(n6715)
         );
  OAI22_X1 U3542 ( .A1(n3100), .A2(n3488), .B1(n7190), .B2(n388), .ZN(n6716)
         );
  OAI22_X1 U3543 ( .A1(n3091), .A2(n3488), .B1(n7190), .B2(n387), .ZN(n6717)
         );
  OAI22_X1 U3544 ( .A1(n3084), .A2(n3488), .B1(n7190), .B2(n386), .ZN(n6718)
         );
  OAI22_X1 U3545 ( .A1(n3075), .A2(n3488), .B1(n7190), .B2(n385), .ZN(n6719)
         );
  OAI22_X1 U3546 ( .A1(n3137), .A2(n3490), .B1(n3306), .B2(n384), .ZN(n6720)
         );
  OAI22_X1 U3547 ( .A1(n3133), .A2(n3490), .B1(n3306), .B2(n383), .ZN(n6721)
         );
  OAI22_X1 U3548 ( .A1(n3118), .A2(n3490), .B1(n3306), .B2(n382), .ZN(n6722)
         );
  OAI22_X1 U3549 ( .A1(n3111), .A2(n3490), .B1(n3306), .B2(n381), .ZN(n6723)
         );
  OAI22_X1 U3550 ( .A1(n3102), .A2(n3490), .B1(n3306), .B2(n380), .ZN(n6724)
         );
  OAI22_X1 U3551 ( .A1(n3093), .A2(n3490), .B1(n3306), .B2(n379), .ZN(n6725)
         );
  OAI22_X1 U3552 ( .A1(n3084), .A2(n3490), .B1(n3306), .B2(n378), .ZN(n6726)
         );
  OAI22_X1 U3553 ( .A1(n3075), .A2(n3490), .B1(n3306), .B2(n377), .ZN(n6727)
         );
  OAI22_X1 U3554 ( .A1(n3137), .A2(n3492), .B1(n7126), .B2(n376), .ZN(n6728)
         );
  OAI22_X1 U3555 ( .A1(n3130), .A2(n3492), .B1(n7126), .B2(n375), .ZN(n6729)
         );
  OAI22_X1 U3556 ( .A1(n7256), .A2(n3492), .B1(n7126), .B2(n374), .ZN(n6730)
         );
  OAI22_X1 U3557 ( .A1(n3111), .A2(n3492), .B1(n7126), .B2(n373), .ZN(n6731)
         );
  OAI22_X1 U3558 ( .A1(n3100), .A2(n3492), .B1(n7126), .B2(n372), .ZN(n6732)
         );
  OAI22_X1 U3559 ( .A1(n3099), .A2(n3492), .B1(n7126), .B2(n371), .ZN(n6733)
         );
  OAI22_X1 U3560 ( .A1(n3084), .A2(n3492), .B1(n7126), .B2(n370), .ZN(n6734)
         );
  OAI22_X1 U3561 ( .A1(n3075), .A2(n3492), .B1(n7126), .B2(n369), .ZN(n6735)
         );
  OAI22_X1 U3562 ( .A1(n3145), .A2(n3493), .B1(n3289), .B2(n368), .ZN(n6736)
         );
  OAI22_X1 U3563 ( .A1(n3132), .A2(n3493), .B1(n3289), .B2(n367), .ZN(n6737)
         );
  OAI22_X1 U3564 ( .A1(n3124), .A2(n3493), .B1(n3289), .B2(n366), .ZN(n6738)
         );
  OAI22_X1 U3565 ( .A1(n3111), .A2(n3493), .B1(n3289), .B2(n365), .ZN(n6739)
         );
  OAI22_X1 U3566 ( .A1(n3103), .A2(n3493), .B1(n3289), .B2(n364), .ZN(n6740)
         );
  OAI22_X1 U3567 ( .A1(n3094), .A2(n3493), .B1(n3289), .B2(n363), .ZN(n6741)
         );
  OAI22_X1 U3568 ( .A1(n3084), .A2(n3493), .B1(n3289), .B2(n362), .ZN(n6742)
         );
  OAI22_X1 U3569 ( .A1(n3075), .A2(n3493), .B1(n3289), .B2(n361), .ZN(n6743)
         );
  OAI22_X1 U3570 ( .A1(n3144), .A2(n3494), .B1(n7237), .B2(n360), .ZN(n6744)
         );
  OAI22_X1 U3571 ( .A1(n3130), .A2(n3494), .B1(n7237), .B2(n359), .ZN(n6745)
         );
  OAI22_X1 U3572 ( .A1(n3127), .A2(n3494), .B1(n7237), .B2(n358), .ZN(n6746)
         );
  OAI22_X1 U3573 ( .A1(n3111), .A2(n3494), .B1(n7237), .B2(n357), .ZN(n6747)
         );
  OAI22_X1 U3574 ( .A1(n3100), .A2(n3494), .B1(n7237), .B2(n356), .ZN(n6748)
         );
  OAI22_X1 U3575 ( .A1(n3098), .A2(n3494), .B1(n7237), .B2(n355), .ZN(n6749)
         );
  OAI22_X1 U3576 ( .A1(n3084), .A2(n3494), .B1(n7237), .B2(n354), .ZN(n6750)
         );
  OAI22_X1 U3577 ( .A1(n3075), .A2(n3494), .B1(n7237), .B2(n353), .ZN(n6751)
         );
  OAI22_X1 U3578 ( .A1(n3143), .A2(n3495), .B1(n7108), .B2(n352), .ZN(n6752)
         );
  OAI22_X1 U3579 ( .A1(n3131), .A2(n3495), .B1(n7108), .B2(n351), .ZN(n6753)
         );
  OAI22_X1 U3580 ( .A1(n3127), .A2(n3495), .B1(n7108), .B2(n350), .ZN(n6754)
         );
  OAI22_X1 U3581 ( .A1(n3111), .A2(n3495), .B1(n7108), .B2(n349), .ZN(n6755)
         );
  OAI22_X1 U3582 ( .A1(n3102), .A2(n3495), .B1(n7108), .B2(n348), .ZN(n6756)
         );
  OAI22_X1 U3583 ( .A1(n3091), .A2(n3495), .B1(n7108), .B2(n347), .ZN(n6757)
         );
  OAI22_X1 U3584 ( .A1(n3084), .A2(n3495), .B1(n7108), .B2(n346), .ZN(n6758)
         );
  OAI22_X1 U3585 ( .A1(n3075), .A2(n3495), .B1(n7108), .B2(n345), .ZN(n6759)
         );
  OAI22_X1 U3586 ( .A1(n3145), .A2(n3496), .B1(n7173), .B2(n344), .ZN(n6760)
         );
  OAI22_X1 U3587 ( .A1(n3130), .A2(n3496), .B1(n7173), .B2(n343), .ZN(n6761)
         );
  OAI22_X1 U3588 ( .A1(n7256), .A2(n3496), .B1(n7173), .B2(n342), .ZN(n6762)
         );
  OAI22_X1 U3589 ( .A1(n3111), .A2(n3496), .B1(n7173), .B2(n341), .ZN(n6763)
         );
  OAI22_X1 U3590 ( .A1(n3100), .A2(n3496), .B1(n7173), .B2(n340), .ZN(n6764)
         );
  OAI22_X1 U3591 ( .A1(n3097), .A2(n3496), .B1(n7173), .B2(n339), .ZN(n6765)
         );
  OAI22_X1 U3592 ( .A1(n3084), .A2(n3496), .B1(n7173), .B2(n338), .ZN(n6766)
         );
  OAI22_X1 U3593 ( .A1(n3075), .A2(n3496), .B1(n7173), .B2(n337), .ZN(n6767)
         );
  OAI22_X1 U3594 ( .A1(n7258), .A2(n3497), .B1(n3273), .B2(n336), .ZN(n6768)
         );
  OAI22_X1 U3595 ( .A1(n3130), .A2(n3497), .B1(n3273), .B2(n335), .ZN(n6769)
         );
  OAI22_X1 U3596 ( .A1(n7256), .A2(n3497), .B1(n3273), .B2(n334), .ZN(n6770)
         );
  OAI22_X1 U3597 ( .A1(n3113), .A2(n3497), .B1(n3273), .B2(n333), .ZN(n6771)
         );
  OAI22_X1 U3598 ( .A1(n3103), .A2(n3497), .B1(n3273), .B2(n332), .ZN(n6772)
         );
  OAI22_X1 U3599 ( .A1(n3093), .A2(n3497), .B1(n3273), .B2(n331), .ZN(n6773)
         );
  OAI22_X1 U3600 ( .A1(n3090), .A2(n3497), .B1(n3273), .B2(n330), .ZN(n6774)
         );
  OAI22_X1 U3601 ( .A1(n3081), .A2(n3497), .B1(n3273), .B2(n329), .ZN(n6775)
         );
  OAI22_X1 U3602 ( .A1(n3137), .A2(n3498), .B1(n7221), .B2(n328), .ZN(n6776)
         );
  OAI22_X1 U3603 ( .A1(n3128), .A2(n3498), .B1(n7221), .B2(n327), .ZN(n6777)
         );
  OAI22_X1 U3604 ( .A1(n7256), .A2(n3498), .B1(n7221), .B2(n326), .ZN(n6778)
         );
  OAI22_X1 U3605 ( .A1(n3113), .A2(n3498), .B1(n7221), .B2(n325), .ZN(n6779)
         );
  OAI22_X1 U3606 ( .A1(n3102), .A2(n3498), .B1(n7221), .B2(n324), .ZN(n6780)
         );
  OAI22_X1 U3607 ( .A1(n3093), .A2(n3498), .B1(n7221), .B2(n323), .ZN(n6781)
         );
  OAI22_X1 U3608 ( .A1(n3083), .A2(n3498), .B1(n7221), .B2(n322), .ZN(n6782)
         );
  OAI22_X1 U3609 ( .A1(n3074), .A2(n3498), .B1(n7221), .B2(n321), .ZN(n6783)
         );
  OAI22_X1 U3610 ( .A1(n3137), .A2(n3499), .B1(n3337), .B2(n320), .ZN(n6784)
         );
  OAI22_X1 U3611 ( .A1(n3129), .A2(n3499), .B1(n3337), .B2(n319), .ZN(n6785)
         );
  OAI22_X1 U3612 ( .A1(n7256), .A2(n3499), .B1(n3337), .B2(n318), .ZN(n6786)
         );
  OAI22_X1 U3613 ( .A1(n3114), .A2(n3499), .B1(n3337), .B2(n317), .ZN(n6787)
         );
  OAI22_X1 U3614 ( .A1(n3103), .A2(n3499), .B1(n3337), .B2(n316), .ZN(n6788)
         );
  OAI22_X1 U3615 ( .A1(n3093), .A2(n3499), .B1(n3337), .B2(n315), .ZN(n6789)
         );
  OAI22_X1 U3616 ( .A1(n3086), .A2(n3499), .B1(n3337), .B2(n314), .ZN(n6790)
         );
  OAI22_X1 U3617 ( .A1(n3077), .A2(n3499), .B1(n3337), .B2(n313), .ZN(n6791)
         );
  OAI22_X1 U3618 ( .A1(n7258), .A2(n3500), .B1(n7157), .B2(n312), .ZN(n6792)
         );
  OAI22_X1 U3619 ( .A1(n3132), .A2(n3500), .B1(n7157), .B2(n311), .ZN(n6793)
         );
  OAI22_X1 U3620 ( .A1(n7256), .A2(n3500), .B1(n7157), .B2(n310), .ZN(n6794)
         );
  OAI22_X1 U3621 ( .A1(n3115), .A2(n3500), .B1(n7157), .B2(n309), .ZN(n6795)
         );
  OAI22_X1 U3622 ( .A1(n3100), .A2(n3500), .B1(n7157), .B2(n308), .ZN(n6796)
         );
  OAI22_X1 U3623 ( .A1(n3093), .A2(n3500), .B1(n7157), .B2(n307), .ZN(n6797)
         );
  OAI22_X1 U3624 ( .A1(n3087), .A2(n3500), .B1(n7157), .B2(n306), .ZN(n6798)
         );
  OAI22_X1 U3625 ( .A1(n3078), .A2(n3500), .B1(n7157), .B2(n305), .ZN(n6799)
         );
  OAI22_X1 U3626 ( .A1(n3143), .A2(n3501), .B1(n3257), .B2(n304), .ZN(n6800)
         );
  OAI22_X1 U3627 ( .A1(n3130), .A2(n3501), .B1(n3257), .B2(n303), .ZN(n6801)
         );
  OAI22_X1 U3628 ( .A1(n3120), .A2(n3501), .B1(n3257), .B2(n302), .ZN(n6802)
         );
  OAI22_X1 U3629 ( .A1(n3112), .A2(n3501), .B1(n3257), .B2(n301), .ZN(n6803)
         );
  OAI22_X1 U3630 ( .A1(n3102), .A2(n3501), .B1(n3257), .B2(n300), .ZN(n6804)
         );
  OAI22_X1 U3631 ( .A1(n3093), .A2(n3501), .B1(n3257), .B2(n299), .ZN(n6805)
         );
  OAI22_X1 U3632 ( .A1(n3088), .A2(n3501), .B1(n3257), .B2(n298), .ZN(n6806)
         );
  OAI22_X1 U3633 ( .A1(n3079), .A2(n3501), .B1(n3257), .B2(n297), .ZN(n6807)
         );
  OAI22_X1 U3634 ( .A1(n3141), .A2(n3502), .B1(n7205), .B2(n296), .ZN(n6808)
         );
  OAI22_X1 U3635 ( .A1(n3128), .A2(n3502), .B1(n7205), .B2(n295), .ZN(n6809)
         );
  OAI22_X1 U3636 ( .A1(n7256), .A2(n3502), .B1(n7205), .B2(n294), .ZN(n6810)
         );
  OAI22_X1 U3637 ( .A1(n3113), .A2(n3502), .B1(n7205), .B2(n293), .ZN(n6811)
         );
  OAI22_X1 U3638 ( .A1(n3100), .A2(n3502), .B1(n7205), .B2(n292), .ZN(n6812)
         );
  OAI22_X1 U3639 ( .A1(n3093), .A2(n3502), .B1(n7205), .B2(n291), .ZN(n6813)
         );
  OAI22_X1 U3640 ( .A1(n3089), .A2(n3502), .B1(n7205), .B2(n290), .ZN(n6814)
         );
  OAI22_X1 U3641 ( .A1(n3080), .A2(n3502), .B1(n7205), .B2(n289), .ZN(n6815)
         );
  OAI22_X1 U3642 ( .A1(n3138), .A2(n3503), .B1(n3321), .B2(n288), .ZN(n6816)
         );
  OAI22_X1 U3643 ( .A1(n3129), .A2(n3503), .B1(n3321), .B2(n287), .ZN(n6817)
         );
  OAI22_X1 U3644 ( .A1(n7256), .A2(n3503), .B1(n3321), .B2(n286), .ZN(n6818)
         );
  OAI22_X1 U3645 ( .A1(n3112), .A2(n3503), .B1(n3321), .B2(n285), .ZN(n6819)
         );
  OAI22_X1 U3646 ( .A1(n3103), .A2(n3503), .B1(n3321), .B2(n284), .ZN(n6820)
         );
  OAI22_X1 U3647 ( .A1(n3093), .A2(n3503), .B1(n3321), .B2(n283), .ZN(n6821)
         );
  OAI22_X1 U3648 ( .A1(n3085), .A2(n3503), .B1(n3321), .B2(n282), .ZN(n6822)
         );
  OAI22_X1 U3649 ( .A1(n3076), .A2(n3503), .B1(n3321), .B2(n281), .ZN(n6823)
         );
  OAI22_X1 U3650 ( .A1(n7258), .A2(n3504), .B1(n7141), .B2(n280), .ZN(n6824)
         );
  OAI22_X1 U3651 ( .A1(n3128), .A2(n3504), .B1(n7141), .B2(n279), .ZN(n6825)
         );
  OAI22_X1 U3652 ( .A1(n7256), .A2(n3504), .B1(n7141), .B2(n278), .ZN(n6826)
         );
  OAI22_X1 U3653 ( .A1(n3114), .A2(n3504), .B1(n7141), .B2(n277), .ZN(n6827)
         );
  OAI22_X1 U3654 ( .A1(n3100), .A2(n3504), .B1(n7141), .B2(n276), .ZN(n6828)
         );
  OAI22_X1 U3655 ( .A1(n3093), .A2(n3504), .B1(n7141), .B2(n275), .ZN(n6829)
         );
  OAI22_X1 U3656 ( .A1(n3086), .A2(n3504), .B1(n7141), .B2(n274), .ZN(n6830)
         );
  OAI22_X1 U3657 ( .A1(n3077), .A2(n3504), .B1(n7141), .B2(n273), .ZN(n6831)
         );
  OAI22_X1 U3658 ( .A1(n7258), .A2(n3505), .B1(n3241), .B2(n272), .ZN(n6832)
         );
  OAI22_X1 U3659 ( .A1(n3129), .A2(n3505), .B1(n3241), .B2(n271), .ZN(n6833)
         );
  OAI22_X1 U3660 ( .A1(n7256), .A2(n3505), .B1(n3241), .B2(n270), .ZN(n6834)
         );
  OAI22_X1 U3661 ( .A1(n3115), .A2(n3505), .B1(n3241), .B2(n269), .ZN(n6835)
         );
  OAI22_X1 U3662 ( .A1(n3102), .A2(n3505), .B1(n3241), .B2(n268), .ZN(n6836)
         );
  OAI22_X1 U3663 ( .A1(n3093), .A2(n3505), .B1(n3241), .B2(n267), .ZN(n6837)
         );
  OAI22_X1 U3664 ( .A1(n3087), .A2(n3505), .B1(n3241), .B2(n266), .ZN(n6838)
         );
  OAI22_X1 U3665 ( .A1(n3078), .A2(n3505), .B1(n3241), .B2(n265), .ZN(n6839)
         );
  OAI22_X1 U3666 ( .A1(n7258), .A2(n3506), .B1(n7189), .B2(n264), .ZN(n6840)
         );
  OAI22_X1 U3667 ( .A1(n3128), .A2(n3506), .B1(n7189), .B2(n263), .ZN(n6841)
         );
  OAI22_X1 U3668 ( .A1(n7256), .A2(n3506), .B1(n7189), .B2(n262), .ZN(n6842)
         );
  OAI22_X1 U3669 ( .A1(n3112), .A2(n3506), .B1(n7189), .B2(n261), .ZN(n6843)
         );
  OAI22_X1 U3670 ( .A1(n3100), .A2(n3506), .B1(n7189), .B2(n260), .ZN(n6844)
         );
  OAI22_X1 U3671 ( .A1(n3093), .A2(n3506), .B1(n7189), .B2(n259), .ZN(n6845)
         );
  OAI22_X1 U3672 ( .A1(n3088), .A2(n3506), .B1(n7189), .B2(n258), .ZN(n6846)
         );
  OAI22_X1 U3673 ( .A1(n3079), .A2(n3506), .B1(n7189), .B2(n257), .ZN(n6847)
         );
  OAI22_X1 U3674 ( .A1(n3139), .A2(n3507), .B1(n3305), .B2(n256), .ZN(n6848)
         );
  OAI22_X1 U3675 ( .A1(n3128), .A2(n3507), .B1(n3305), .B2(n255), .ZN(n6849)
         );
  OAI22_X1 U3676 ( .A1(n3121), .A2(n3507), .B1(n3305), .B2(n254), .ZN(n6850)
         );
  OAI22_X1 U3677 ( .A1(n3113), .A2(n3507), .B1(n3305), .B2(n253), .ZN(n6851)
         );
  OAI22_X1 U3678 ( .A1(n3103), .A2(n3507), .B1(n3305), .B2(n252), .ZN(n6852)
         );
  OAI22_X1 U3679 ( .A1(n3093), .A2(n3507), .B1(n3305), .B2(n251), .ZN(n6853)
         );
  OAI22_X1 U3680 ( .A1(n3089), .A2(n3507), .B1(n3305), .B2(n250), .ZN(n6854)
         );
  OAI22_X1 U3681 ( .A1(n3080), .A2(n3507), .B1(n3305), .B2(n249), .ZN(n6855)
         );
  OAI22_X1 U3682 ( .A1(n3145), .A2(n3509), .B1(n7125), .B2(n248), .ZN(n6856)
         );
  OAI22_X1 U3683 ( .A1(n3136), .A2(n3509), .B1(n7125), .B2(n247), .ZN(n6857)
         );
  OAI22_X1 U3684 ( .A1(n3127), .A2(n3509), .B1(n7125), .B2(n246), .ZN(n6858)
         );
  OAI22_X1 U3685 ( .A1(n3115), .A2(n3509), .B1(n7125), .B2(n245), .ZN(n6859)
         );
  OAI22_X1 U3686 ( .A1(n3100), .A2(n3509), .B1(n7125), .B2(n244), .ZN(n6860)
         );
  OAI22_X1 U3687 ( .A1(n3093), .A2(n3509), .B1(n7125), .B2(n243), .ZN(n6861)
         );
  OAI22_X1 U3688 ( .A1(n3085), .A2(n3509), .B1(n7125), .B2(n242), .ZN(n6862)
         );
  OAI22_X1 U3689 ( .A1(n3076), .A2(n3509), .B1(n7125), .B2(n241), .ZN(n6863)
         );
  OAI22_X1 U3690 ( .A1(n3145), .A2(n3510), .B1(n3288), .B2(n240), .ZN(n6864)
         );
  OAI22_X1 U3691 ( .A1(n3136), .A2(n3510), .B1(n3288), .B2(n239), .ZN(n6865)
         );
  OAI22_X1 U3692 ( .A1(n3127), .A2(n3510), .B1(n3288), .B2(n238), .ZN(n6866)
         );
  OAI22_X1 U3693 ( .A1(n3114), .A2(n3510), .B1(n3288), .B2(n237), .ZN(n6867)
         );
  OAI22_X1 U3694 ( .A1(n3104), .A2(n3510), .B1(n3288), .B2(n236), .ZN(n6868)
         );
  OAI22_X1 U3695 ( .A1(n3093), .A2(n3510), .B1(n3288), .B2(n235), .ZN(n6869)
         );
  OAI22_X1 U3696 ( .A1(n3086), .A2(n3510), .B1(n3288), .B2(n234), .ZN(n6870)
         );
  OAI22_X1 U3697 ( .A1(n3077), .A2(n3510), .B1(n3288), .B2(n233), .ZN(n6871)
         );
  OAI22_X1 U3698 ( .A1(n3145), .A2(n3511), .B1(n7236), .B2(n232), .ZN(n6872)
         );
  OAI22_X1 U3699 ( .A1(n3136), .A2(n3511), .B1(n7236), .B2(n231), .ZN(n6873)
         );
  OAI22_X1 U3700 ( .A1(n3127), .A2(n3511), .B1(n7236), .B2(n230), .ZN(n6874)
         );
  OAI22_X1 U3701 ( .A1(n3112), .A2(n3511), .B1(n7236), .B2(n229), .ZN(n6875)
         );
  OAI22_X1 U3702 ( .A1(n3101), .A2(n3511), .B1(n7236), .B2(n228), .ZN(n6876)
         );
  OAI22_X1 U3703 ( .A1(n3094), .A2(n3511), .B1(n7236), .B2(n227), .ZN(n6877)
         );
  OAI22_X1 U3704 ( .A1(n3085), .A2(n3511), .B1(n7236), .B2(n226), .ZN(n6878)
         );
  OAI22_X1 U3705 ( .A1(n3076), .A2(n3511), .B1(n7236), .B2(n225), .ZN(n6879)
         );
  OAI22_X1 U3706 ( .A1(n3145), .A2(n3512), .B1(n7107), .B2(n224), .ZN(n6880)
         );
  OAI22_X1 U3707 ( .A1(n3136), .A2(n3512), .B1(n7107), .B2(n223), .ZN(n6881)
         );
  OAI22_X1 U3708 ( .A1(n3127), .A2(n3512), .B1(n7107), .B2(n222), .ZN(n6882)
         );
  OAI22_X1 U3709 ( .A1(n3112), .A2(n3512), .B1(n7107), .B2(n221), .ZN(n6883)
         );
  OAI22_X1 U3710 ( .A1(n3101), .A2(n3512), .B1(n7107), .B2(n220), .ZN(n6884)
         );
  OAI22_X1 U3711 ( .A1(n3094), .A2(n3512), .B1(n7107), .B2(n219), .ZN(n6885)
         );
  OAI22_X1 U3712 ( .A1(n3085), .A2(n3512), .B1(n7107), .B2(n218), .ZN(n6886)
         );
  OAI22_X1 U3713 ( .A1(n3076), .A2(n3512), .B1(n7107), .B2(n217), .ZN(n6887)
         );
  OAI22_X1 U3714 ( .A1(n3145), .A2(n3513), .B1(n7172), .B2(n216), .ZN(n6888)
         );
  OAI22_X1 U3715 ( .A1(n3136), .A2(n3513), .B1(n7172), .B2(n215), .ZN(n6889)
         );
  OAI22_X1 U3716 ( .A1(n3127), .A2(n3513), .B1(n7172), .B2(n214), .ZN(n6890)
         );
  OAI22_X1 U3717 ( .A1(n3112), .A2(n3513), .B1(n7172), .B2(n213), .ZN(n6891)
         );
  OAI22_X1 U3718 ( .A1(n3101), .A2(n3513), .B1(n7172), .B2(n212), .ZN(n6892)
         );
  OAI22_X1 U3719 ( .A1(n3094), .A2(n3513), .B1(n7172), .B2(n211), .ZN(n6893)
         );
  OAI22_X1 U3720 ( .A1(n3085), .A2(n3513), .B1(n7172), .B2(n210), .ZN(n6894)
         );
  OAI22_X1 U3721 ( .A1(n3076), .A2(n3513), .B1(n7172), .B2(n209), .ZN(n6895)
         );
  OAI22_X1 U3722 ( .A1(n3145), .A2(n3514), .B1(n3272), .B2(n208), .ZN(n6896)
         );
  OAI22_X1 U3723 ( .A1(n3136), .A2(n3514), .B1(n3272), .B2(n207), .ZN(n6897)
         );
  OAI22_X1 U3724 ( .A1(n3127), .A2(n3514), .B1(n3272), .B2(n206), .ZN(n6898)
         );
  OAI22_X1 U3725 ( .A1(n3112), .A2(n3514), .B1(n3272), .B2(n205), .ZN(n6899)
         );
  OAI22_X1 U3726 ( .A1(n3101), .A2(n3514), .B1(n3272), .B2(n204), .ZN(n6900)
         );
  OAI22_X1 U3727 ( .A1(n3094), .A2(n3514), .B1(n3272), .B2(n203), .ZN(n6901)
         );
  OAI22_X1 U3728 ( .A1(n3085), .A2(n3514), .B1(n3272), .B2(n202), .ZN(n6902)
         );
  OAI22_X1 U3729 ( .A1(n3076), .A2(n3514), .B1(n3272), .B2(n201), .ZN(n6903)
         );
  OAI22_X1 U3730 ( .A1(n3145), .A2(n3515), .B1(n7220), .B2(n200), .ZN(n6904)
         );
  OAI22_X1 U3731 ( .A1(n3136), .A2(n3515), .B1(n7220), .B2(n199), .ZN(n6905)
         );
  OAI22_X1 U3732 ( .A1(n3127), .A2(n3515), .B1(n7220), .B2(n198), .ZN(n6906)
         );
  OAI22_X1 U3733 ( .A1(n3112), .A2(n3515), .B1(n7220), .B2(n197), .ZN(n6907)
         );
  OAI22_X1 U3734 ( .A1(n3101), .A2(n3515), .B1(n7220), .B2(n196), .ZN(n6908)
         );
  OAI22_X1 U3735 ( .A1(n3094), .A2(n3515), .B1(n7220), .B2(n195), .ZN(n6909)
         );
  OAI22_X1 U3736 ( .A1(n3085), .A2(n3515), .B1(n7220), .B2(n194), .ZN(n6910)
         );
  OAI22_X1 U3737 ( .A1(n3076), .A2(n3515), .B1(n7220), .B2(n193), .ZN(n6911)
         );
  OAI22_X1 U3738 ( .A1(n3145), .A2(n3516), .B1(n3336), .B2(n192), .ZN(n6912)
         );
  OAI22_X1 U3739 ( .A1(n3136), .A2(n3516), .B1(n3336), .B2(n191), .ZN(n6913)
         );
  OAI22_X1 U3740 ( .A1(n3127), .A2(n3516), .B1(n3336), .B2(n190), .ZN(n6914)
         );
  OAI22_X1 U3741 ( .A1(n3112), .A2(n3516), .B1(n3336), .B2(n189), .ZN(n6915)
         );
  OAI22_X1 U3742 ( .A1(n3101), .A2(n3516), .B1(n3336), .B2(n188), .ZN(n6916)
         );
  OAI22_X1 U3743 ( .A1(n3094), .A2(n3516), .B1(n3336), .B2(n187), .ZN(n6917)
         );
  OAI22_X1 U3744 ( .A1(n3085), .A2(n3516), .B1(n3336), .B2(n186), .ZN(n6918)
         );
  OAI22_X1 U3745 ( .A1(n3076), .A2(n3516), .B1(n3336), .B2(n185), .ZN(n6919)
         );
  OAI22_X1 U3746 ( .A1(n3145), .A2(n3517), .B1(n7156), .B2(n184), .ZN(n6920)
         );
  OAI22_X1 U3747 ( .A1(n3136), .A2(n3517), .B1(n7156), .B2(n183), .ZN(n6921)
         );
  OAI22_X1 U3748 ( .A1(n3127), .A2(n3517), .B1(n7156), .B2(n182), .ZN(n6922)
         );
  OAI22_X1 U3749 ( .A1(n3112), .A2(n3517), .B1(n7156), .B2(n181), .ZN(n6923)
         );
  OAI22_X1 U3750 ( .A1(n3101), .A2(n3517), .B1(n7156), .B2(n180), .ZN(n6924)
         );
  OAI22_X1 U3751 ( .A1(n3094), .A2(n3517), .B1(n7156), .B2(n179), .ZN(n6925)
         );
  OAI22_X1 U3752 ( .A1(n3085), .A2(n3517), .B1(n7156), .B2(n178), .ZN(n6926)
         );
  OAI22_X1 U3753 ( .A1(n3076), .A2(n3517), .B1(n7156), .B2(n177), .ZN(n6927)
         );
  OAI22_X1 U3754 ( .A1(n3144), .A2(n3518), .B1(n3256), .B2(n176), .ZN(n6928)
         );
  OAI22_X1 U3755 ( .A1(n3135), .A2(n3518), .B1(n3256), .B2(n175), .ZN(n6929)
         );
  OAI22_X1 U3756 ( .A1(n3126), .A2(n3518), .B1(n3256), .B2(n174), .ZN(n6930)
         );
  OAI22_X1 U3757 ( .A1(n3112), .A2(n3518), .B1(n3256), .B2(n173), .ZN(n6931)
         );
  OAI22_X1 U3758 ( .A1(n3101), .A2(n3518), .B1(n3256), .B2(n172), .ZN(n6932)
         );
  OAI22_X1 U3759 ( .A1(n3094), .A2(n3518), .B1(n3256), .B2(n171), .ZN(n6933)
         );
  OAI22_X1 U3760 ( .A1(n3085), .A2(n3518), .B1(n3256), .B2(n170), .ZN(n6934)
         );
  OAI22_X1 U3761 ( .A1(n3076), .A2(n3518), .B1(n3256), .B2(n169), .ZN(n6935)
         );
  OAI22_X1 U3762 ( .A1(n3144), .A2(n3519), .B1(n7204), .B2(n168), .ZN(n6936)
         );
  OAI22_X1 U3763 ( .A1(n3136), .A2(n3519), .B1(n7204), .B2(n167), .ZN(n6937)
         );
  OAI22_X1 U3764 ( .A1(n3126), .A2(n3519), .B1(n7204), .B2(n166), .ZN(n6938)
         );
  OAI22_X1 U3765 ( .A1(n3112), .A2(n3519), .B1(n7204), .B2(n165), .ZN(n6939)
         );
  OAI22_X1 U3766 ( .A1(n3101), .A2(n3519), .B1(n7204), .B2(n164), .ZN(n6940)
         );
  OAI22_X1 U3767 ( .A1(n3094), .A2(n3519), .B1(n7204), .B2(n163), .ZN(n6941)
         );
  OAI22_X1 U3768 ( .A1(n3085), .A2(n3519), .B1(n7204), .B2(n162), .ZN(n6942)
         );
  OAI22_X1 U3769 ( .A1(n3076), .A2(n3519), .B1(n7204), .B2(n161), .ZN(n6943)
         );
  OAI22_X1 U3770 ( .A1(n3144), .A2(n3520), .B1(n3320), .B2(n160), .ZN(n6944)
         );
  OAI22_X1 U3771 ( .A1(n3134), .A2(n3520), .B1(n3320), .B2(n159), .ZN(n6945)
         );
  OAI22_X1 U3772 ( .A1(n3126), .A2(n3520), .B1(n3320), .B2(n158), .ZN(n6946)
         );
  OAI22_X1 U3773 ( .A1(n3112), .A2(n3520), .B1(n3320), .B2(n157), .ZN(n6947)
         );
  OAI22_X1 U3774 ( .A1(n3101), .A2(n3520), .B1(n3320), .B2(n156), .ZN(n6948)
         );
  OAI22_X1 U3775 ( .A1(n3094), .A2(n3520), .B1(n3320), .B2(n155), .ZN(n6949)
         );
  OAI22_X1 U3776 ( .A1(n3085), .A2(n3520), .B1(n3320), .B2(n154), .ZN(n6950)
         );
  OAI22_X1 U3777 ( .A1(n3076), .A2(n3520), .B1(n3320), .B2(n153), .ZN(n6951)
         );
  OAI22_X1 U3778 ( .A1(n3144), .A2(n3521), .B1(n7140), .B2(n152), .ZN(n6952)
         );
  OAI22_X1 U3779 ( .A1(n3133), .A2(n3521), .B1(n7140), .B2(n151), .ZN(n6953)
         );
  OAI22_X1 U3780 ( .A1(n3126), .A2(n3521), .B1(n7140), .B2(n150), .ZN(n6954)
         );
  OAI22_X1 U3781 ( .A1(n3112), .A2(n3521), .B1(n7140), .B2(n149), .ZN(n6955)
         );
  OAI22_X1 U3782 ( .A1(n3101), .A2(n3521), .B1(n7140), .B2(n148), .ZN(n6956)
         );
  OAI22_X1 U3783 ( .A1(n3094), .A2(n3521), .B1(n7140), .B2(n147), .ZN(n6957)
         );
  OAI22_X1 U3784 ( .A1(n3085), .A2(n3521), .B1(n7140), .B2(n146), .ZN(n6958)
         );
  OAI22_X1 U3785 ( .A1(n3076), .A2(n3521), .B1(n7140), .B2(n145), .ZN(n6959)
         );
  OAI22_X1 U3786 ( .A1(n3144), .A2(n3522), .B1(n3240), .B2(n144), .ZN(n6960)
         );
  OAI22_X1 U3787 ( .A1(n3132), .A2(n3522), .B1(n3240), .B2(n143), .ZN(n6961)
         );
  OAI22_X1 U3788 ( .A1(n3126), .A2(n3522), .B1(n3240), .B2(n142), .ZN(n6962)
         );
  OAI22_X1 U3789 ( .A1(n3112), .A2(n3522), .B1(n3240), .B2(n141), .ZN(n6963)
         );
  OAI22_X1 U3790 ( .A1(n3101), .A2(n3522), .B1(n3240), .B2(n140), .ZN(n6964)
         );
  OAI22_X1 U3791 ( .A1(n3094), .A2(n3522), .B1(n3240), .B2(n139), .ZN(n6965)
         );
  OAI22_X1 U3792 ( .A1(n3085), .A2(n3522), .B1(n3240), .B2(n138), .ZN(n6966)
         );
  OAI22_X1 U3793 ( .A1(n3076), .A2(n3522), .B1(n3240), .B2(n137), .ZN(n6967)
         );
  OAI22_X1 U3794 ( .A1(n3144), .A2(n3523), .B1(n7188), .B2(n136), .ZN(n6968)
         );
  OAI22_X1 U3795 ( .A1(n3131), .A2(n3523), .B1(n7188), .B2(n135), .ZN(n6969)
         );
  OAI22_X1 U3796 ( .A1(n3126), .A2(n3523), .B1(n7188), .B2(n134), .ZN(n6970)
         );
  OAI22_X1 U3797 ( .A1(n3112), .A2(n3523), .B1(n7188), .B2(n133), .ZN(n6971)
         );
  OAI22_X1 U3798 ( .A1(n3101), .A2(n3523), .B1(n7188), .B2(n132), .ZN(n6972)
         );
  OAI22_X1 U3799 ( .A1(n3094), .A2(n3523), .B1(n7188), .B2(n131), .ZN(n6973)
         );
  OAI22_X1 U3800 ( .A1(n3085), .A2(n3523), .B1(n7188), .B2(n130), .ZN(n6974)
         );
  OAI22_X1 U3801 ( .A1(n3076), .A2(n3523), .B1(n7188), .B2(n129), .ZN(n6975)
         );
  OAI22_X1 U3802 ( .A1(n3144), .A2(n3524), .B1(n3304), .B2(n128), .ZN(n6976)
         );
  OAI22_X1 U3803 ( .A1(n3128), .A2(n3524), .B1(n3304), .B2(n127), .ZN(n6977)
         );
  OAI22_X1 U3804 ( .A1(n3126), .A2(n3524), .B1(n3304), .B2(n126), .ZN(n6978)
         );
  OAI22_X1 U3805 ( .A1(n3113), .A2(n3524), .B1(n3304), .B2(n125), .ZN(n6979)
         );
  OAI22_X1 U3806 ( .A1(n3108), .A2(n3524), .B1(n3304), .B2(n124), .ZN(n6980)
         );
  OAI22_X1 U3807 ( .A1(n3095), .A2(n3524), .B1(n3304), .B2(n123), .ZN(n6981)
         );
  OAI22_X1 U3808 ( .A1(n3086), .A2(n3524), .B1(n3304), .B2(n122), .ZN(n6982)
         );
  OAI22_X1 U3809 ( .A1(n3077), .A2(n3524), .B1(n3304), .B2(n121), .ZN(n6983)
         );
  OAI22_X1 U3810 ( .A1(n3144), .A2(n3526), .B1(n7124), .B2(n120), .ZN(n6984)
         );
  OAI22_X1 U3811 ( .A1(n3136), .A2(n3526), .B1(n7124), .B2(n119), .ZN(n6985)
         );
  OAI22_X1 U3812 ( .A1(n3126), .A2(n3526), .B1(n7124), .B2(n118), .ZN(n6986)
         );
  OAI22_X1 U3813 ( .A1(n3113), .A2(n3526), .B1(n7124), .B2(n117), .ZN(n6987)
         );
  OAI22_X1 U3814 ( .A1(n3107), .A2(n3526), .B1(n7124), .B2(n116), .ZN(n6988)
         );
  OAI22_X1 U3815 ( .A1(n3095), .A2(n3526), .B1(n7124), .B2(n115), .ZN(n6989)
         );
  OAI22_X1 U3816 ( .A1(n3086), .A2(n3526), .B1(n7124), .B2(n114), .ZN(n6990)
         );
  OAI22_X1 U3817 ( .A1(n3077), .A2(n3526), .B1(n7124), .B2(n113), .ZN(n6991)
         );
  OAI22_X1 U3818 ( .A1(n3144), .A2(n3527), .B1(n3287), .B2(n112), .ZN(n6992)
         );
  OAI22_X1 U3819 ( .A1(n3133), .A2(n3527), .B1(n3287), .B2(n111), .ZN(n6993)
         );
  OAI22_X1 U3820 ( .A1(n3126), .A2(n3527), .B1(n3287), .B2(n110), .ZN(n6994)
         );
  OAI22_X1 U3821 ( .A1(n3113), .A2(n3527), .B1(n3287), .B2(n109), .ZN(n6995)
         );
  OAI22_X1 U3822 ( .A1(n3108), .A2(n3527), .B1(n3287), .B2(n108), .ZN(n6996)
         );
  OAI22_X1 U3823 ( .A1(n3095), .A2(n3527), .B1(n3287), .B2(n107), .ZN(n6997)
         );
  OAI22_X1 U3824 ( .A1(n3086), .A2(n3527), .B1(n3287), .B2(n106), .ZN(n6998)
         );
  OAI22_X1 U3825 ( .A1(n3077), .A2(n3527), .B1(n3287), .B2(n105), .ZN(n6999)
         );
  OAI22_X1 U3826 ( .A1(n3144), .A2(n3528), .B1(n7235), .B2(n104), .ZN(n7000)
         );
  OAI22_X1 U3827 ( .A1(n3135), .A2(n3528), .B1(n7235), .B2(n103), .ZN(n7001)
         );
  OAI22_X1 U3828 ( .A1(n3126), .A2(n3528), .B1(n7235), .B2(n102), .ZN(n7002)
         );
  OAI22_X1 U3829 ( .A1(n3113), .A2(n3528), .B1(n7235), .B2(n101), .ZN(n7003)
         );
  OAI22_X1 U3830 ( .A1(n3107), .A2(n3528), .B1(n7235), .B2(n100), .ZN(n7004)
         );
  OAI22_X1 U3831 ( .A1(n3095), .A2(n3528), .B1(n7235), .B2(n99), .ZN(n7005) );
  OAI22_X1 U3832 ( .A1(n3086), .A2(n3528), .B1(n7235), .B2(n98), .ZN(n7006) );
  OAI22_X1 U3833 ( .A1(n3077), .A2(n3528), .B1(n7235), .B2(n97), .ZN(n7007) );
  OAI22_X1 U3834 ( .A1(n3144), .A2(n3529), .B1(n7106), .B2(n96), .ZN(n7008) );
  OAI22_X1 U3835 ( .A1(n3136), .A2(n3529), .B1(n7106), .B2(n95), .ZN(n7009) );
  OAI22_X1 U3836 ( .A1(n3126), .A2(n3529), .B1(n7106), .B2(n94), .ZN(n7010) );
  OAI22_X1 U3837 ( .A1(n3113), .A2(n3529), .B1(n7106), .B2(n93), .ZN(n7011) );
  OAI22_X1 U3838 ( .A1(n3108), .A2(n3529), .B1(n7106), .B2(n92), .ZN(n7012) );
  OAI22_X1 U3839 ( .A1(n3095), .A2(n3529), .B1(n7106), .B2(n91), .ZN(n7013) );
  OAI22_X1 U3840 ( .A1(n3086), .A2(n3529), .B1(n7106), .B2(n90), .ZN(n7014) );
  OAI22_X1 U3841 ( .A1(n3077), .A2(n3529), .B1(n7106), .B2(n89), .ZN(n7015) );
  OAI22_X1 U3842 ( .A1(n3144), .A2(n3530), .B1(n7171), .B2(n88), .ZN(n7016) );
  OAI22_X1 U3843 ( .A1(n3134), .A2(n3530), .B1(n7171), .B2(n87), .ZN(n7017) );
  OAI22_X1 U3844 ( .A1(n3126), .A2(n3530), .B1(n7171), .B2(n86), .ZN(n7018) );
  OAI22_X1 U3845 ( .A1(n3113), .A2(n3530), .B1(n7171), .B2(n85), .ZN(n7019) );
  OAI22_X1 U3846 ( .A1(n3107), .A2(n3530), .B1(n7171), .B2(n84), .ZN(n7020) );
  OAI22_X1 U3847 ( .A1(n3095), .A2(n3530), .B1(n7171), .B2(n83), .ZN(n7021) );
  OAI22_X1 U3848 ( .A1(n3086), .A2(n3530), .B1(n7171), .B2(n82), .ZN(n7022) );
  OAI22_X1 U3849 ( .A1(n3077), .A2(n3530), .B1(n7171), .B2(n81), .ZN(n7023) );
  OAI22_X1 U3850 ( .A1(n3144), .A2(n3531), .B1(n3271), .B2(n80), .ZN(n7024) );
  OAI22_X1 U3851 ( .A1(n3133), .A2(n3531), .B1(n3271), .B2(n79), .ZN(n7025) );
  OAI22_X1 U3852 ( .A1(n3126), .A2(n3531), .B1(n3271), .B2(n78), .ZN(n7026) );
  OAI22_X1 U3853 ( .A1(n3113), .A2(n3531), .B1(n3271), .B2(n77), .ZN(n7027) );
  OAI22_X1 U3854 ( .A1(n3108), .A2(n3531), .B1(n3271), .B2(n76), .ZN(n7028) );
  OAI22_X1 U3855 ( .A1(n3095), .A2(n3531), .B1(n3271), .B2(n75), .ZN(n7029) );
  OAI22_X1 U3856 ( .A1(n3086), .A2(n3531), .B1(n3271), .B2(n74), .ZN(n7030) );
  OAI22_X1 U3857 ( .A1(n3077), .A2(n3531), .B1(n3271), .B2(n73), .ZN(n7031) );
  OAI22_X1 U3858 ( .A1(n3143), .A2(n3532), .B1(n7219), .B2(n72), .ZN(n7032) );
  OAI22_X1 U3859 ( .A1(n3135), .A2(n3532), .B1(n7219), .B2(n71), .ZN(n7033) );
  OAI22_X1 U3860 ( .A1(n3125), .A2(n3532), .B1(n7219), .B2(n70), .ZN(n7034) );
  OAI22_X1 U3861 ( .A1(n3113), .A2(n3532), .B1(n7219), .B2(n69), .ZN(n7035) );
  OAI22_X1 U3862 ( .A1(n3107), .A2(n3532), .B1(n7219), .B2(n68), .ZN(n7036) );
  OAI22_X1 U3863 ( .A1(n3095), .A2(n3532), .B1(n7219), .B2(n67), .ZN(n7037) );
  OAI22_X1 U3864 ( .A1(n3086), .A2(n3532), .B1(n7219), .B2(n66), .ZN(n7038) );
  OAI22_X1 U3865 ( .A1(n3077), .A2(n3532), .B1(n7219), .B2(n65), .ZN(n7039) );
  OAI22_X1 U3866 ( .A1(n3143), .A2(n3533), .B1(n3335), .B2(n64), .ZN(n7040) );
  OAI22_X1 U3867 ( .A1(n3135), .A2(n3533), .B1(n3335), .B2(n63), .ZN(n7041) );
  OAI22_X1 U3868 ( .A1(n3125), .A2(n3533), .B1(n3335), .B2(n62), .ZN(n7042) );
  OAI22_X1 U3869 ( .A1(n3113), .A2(n3533), .B1(n3335), .B2(n61), .ZN(n7043) );
  OAI22_X1 U3870 ( .A1(n3108), .A2(n3533), .B1(n3335), .B2(n60), .ZN(n7044) );
  OAI22_X1 U3871 ( .A1(n3095), .A2(n3533), .B1(n3335), .B2(n59), .ZN(n7045) );
  OAI22_X1 U3872 ( .A1(n3086), .A2(n3533), .B1(n3335), .B2(n58), .ZN(n7046) );
  OAI22_X1 U3873 ( .A1(n3077), .A2(n3533), .B1(n3335), .B2(n57), .ZN(n7047) );
  OAI22_X1 U3874 ( .A1(n3143), .A2(n3534), .B1(n7155), .B2(n56), .ZN(n7048) );
  OAI22_X1 U3875 ( .A1(n3135), .A2(n3534), .B1(n7155), .B2(n55), .ZN(n7049) );
  OAI22_X1 U3876 ( .A1(n3125), .A2(n3534), .B1(n7155), .B2(n54), .ZN(n7050) );
  OAI22_X1 U3877 ( .A1(n3113), .A2(n3534), .B1(n7155), .B2(n53), .ZN(n7051) );
  OAI22_X1 U3878 ( .A1(n3107), .A2(n3534), .B1(n7155), .B2(n52), .ZN(n7052) );
  OAI22_X1 U3879 ( .A1(n3095), .A2(n3534), .B1(n7155), .B2(n51), .ZN(n7053) );
  OAI22_X1 U3880 ( .A1(n3086), .A2(n3534), .B1(n7155), .B2(n50), .ZN(n7054) );
  OAI22_X1 U3881 ( .A1(n3077), .A2(n3534), .B1(n7155), .B2(n49), .ZN(n7055) );
  OAI22_X1 U3882 ( .A1(n3143), .A2(n3535), .B1(n3255), .B2(n48), .ZN(n7056) );
  OAI22_X1 U3883 ( .A1(n3135), .A2(n3535), .B1(n3255), .B2(n47), .ZN(n7057) );
  OAI22_X1 U3884 ( .A1(n3125), .A2(n3535), .B1(n3255), .B2(n46), .ZN(n7058) );
  OAI22_X1 U3885 ( .A1(n3113), .A2(n3535), .B1(n3255), .B2(n45), .ZN(n7059) );
  OAI22_X1 U3886 ( .A1(n3108), .A2(n3535), .B1(n3255), .B2(n44), .ZN(n7060) );
  OAI22_X1 U3887 ( .A1(n3095), .A2(n3535), .B1(n3255), .B2(n43), .ZN(n7061) );
  OAI22_X1 U3888 ( .A1(n3086), .A2(n3535), .B1(n3255), .B2(n42), .ZN(n7062) );
  OAI22_X1 U3889 ( .A1(n3077), .A2(n3535), .B1(n3255), .B2(n41), .ZN(n7063) );
  OAI22_X1 U3890 ( .A1(n3143), .A2(n3536), .B1(n7203), .B2(n40), .ZN(n7064) );
  OAI22_X1 U3891 ( .A1(n3135), .A2(n3536), .B1(n7203), .B2(n39), .ZN(n7065) );
  OAI22_X1 U3892 ( .A1(n3125), .A2(n3536), .B1(n7203), .B2(n38), .ZN(n7066) );
  OAI22_X1 U3893 ( .A1(n3113), .A2(n3536), .B1(n7203), .B2(n37), .ZN(n7067) );
  OAI22_X1 U3894 ( .A1(n3107), .A2(n3536), .B1(n7203), .B2(n36), .ZN(n7068) );
  OAI22_X1 U3895 ( .A1(n3095), .A2(n3536), .B1(n7203), .B2(n35), .ZN(n7069) );
  OAI22_X1 U3896 ( .A1(n3086), .A2(n3536), .B1(n7203), .B2(n34), .ZN(n7070) );
  OAI22_X1 U3897 ( .A1(n3077), .A2(n3536), .B1(n7203), .B2(n33), .ZN(n7071) );
  OAI22_X1 U3898 ( .A1(n3143), .A2(n3537), .B1(n3319), .B2(n32), .ZN(n7072) );
  OAI22_X1 U3899 ( .A1(n3135), .A2(n3537), .B1(n3319), .B2(n31), .ZN(n7073) );
  OAI22_X1 U3900 ( .A1(n3125), .A2(n3537), .B1(n3319), .B2(n30), .ZN(n7074) );
  OAI22_X1 U3901 ( .A1(n3113), .A2(n3537), .B1(n3319), .B2(n29), .ZN(n7075) );
  OAI22_X1 U3902 ( .A1(n3108), .A2(n3537), .B1(n3319), .B2(n28), .ZN(n7076) );
  OAI22_X1 U3903 ( .A1(n3095), .A2(n3537), .B1(n3319), .B2(n27), .ZN(n7077) );
  OAI22_X1 U3904 ( .A1(n3086), .A2(n3537), .B1(n3319), .B2(n26), .ZN(n7078) );
  OAI22_X1 U3905 ( .A1(n3077), .A2(n3537), .B1(n3319), .B2(n25), .ZN(n7079) );
  OAI22_X1 U3906 ( .A1(n3143), .A2(n3538), .B1(n7139), .B2(n24), .ZN(n7080) );
  OAI22_X1 U3907 ( .A1(n3135), .A2(n3538), .B1(n7139), .B2(n23), .ZN(n7081) );
  OAI22_X1 U3908 ( .A1(n3125), .A2(n3538), .B1(n7139), .B2(n22), .ZN(n7082) );
  OAI22_X1 U3909 ( .A1(n3114), .A2(n3538), .B1(n7139), .B2(n21), .ZN(n7083) );
  OAI22_X1 U3910 ( .A1(n3102), .A2(n3538), .B1(n7139), .B2(n20), .ZN(n7084) );
  OAI22_X1 U3911 ( .A1(n3096), .A2(n3538), .B1(n7139), .B2(n19), .ZN(n7085) );
  OAI22_X1 U3912 ( .A1(n3087), .A2(n3538), .B1(n7139), .B2(n18), .ZN(n7086) );
  OAI22_X1 U3913 ( .A1(n3078), .A2(n3538), .B1(n7139), .B2(n17), .ZN(n7087) );
  OAI22_X1 U3914 ( .A1(n3143), .A2(n3539), .B1(n3239), .B2(n16), .ZN(n7088) );
  OAI22_X1 U3915 ( .A1(n3135), .A2(n3539), .B1(n3239), .B2(n15), .ZN(n7089) );
  OAI22_X1 U3916 ( .A1(n3125), .A2(n3539), .B1(n3239), .B2(n14), .ZN(n7090) );
  OAI22_X1 U3917 ( .A1(n7255), .A2(n3539), .B1(n3239), .B2(n13), .ZN(n7091) );
  OAI22_X1 U3918 ( .A1(n3102), .A2(n3539), .B1(n3239), .B2(n12), .ZN(n7092) );
  OAI22_X1 U3919 ( .A1(n3096), .A2(n3539), .B1(n3239), .B2(n11), .ZN(n7093) );
  OAI22_X1 U3920 ( .A1(n3087), .A2(n3539), .B1(n3239), .B2(n10), .ZN(n7094) );
  OAI22_X1 U3921 ( .A1(n3078), .A2(n3539), .B1(n3239), .B2(n9), .ZN(n7095) );
  OAI22_X1 U3922 ( .A1(n3143), .A2(n3540), .B1(n7187), .B2(n8), .ZN(n7096) );
  OAI22_X1 U3923 ( .A1(n3135), .A2(n3540), .B1(n7187), .B2(n7), .ZN(n7097) );
  OAI22_X1 U3924 ( .A1(n3125), .A2(n3540), .B1(n7187), .B2(n6), .ZN(n7098) );
  OAI22_X1 U3925 ( .A1(n3109), .A2(n3540), .B1(n7187), .B2(n5), .ZN(n7099) );
  OAI22_X1 U3926 ( .A1(n3102), .A2(n3540), .B1(n7187), .B2(n4), .ZN(n7100) );
  OAI22_X1 U3927 ( .A1(n3096), .A2(n3540), .B1(n7187), .B2(n3), .ZN(n7101) );
  OAI22_X1 U3928 ( .A1(n3087), .A2(n3540), .B1(n7187), .B2(n2), .ZN(n7102) );
  OAI22_X1 U3929 ( .A1(n3078), .A2(n3540), .B1(n7187), .B2(n1), .ZN(n7103) );
  OAI22_X1 U3930 ( .A1(n7255), .A2(n3350), .B1(n3296), .B2(n1949), .ZN(n5843)
         );
  OAI22_X1 U3931 ( .A1(n7254), .A2(n3350), .B1(n3296), .B2(n1948), .ZN(n5844)
         );
  OAI22_X1 U3932 ( .A1(n3091), .A2(n3350), .B1(n3296), .B2(n1947), .ZN(n5845)
         );
  OAI22_X1 U3933 ( .A1(n7252), .A2(n3350), .B1(n3296), .B2(n1946), .ZN(n5846)
         );
  OAI22_X1 U3934 ( .A1(n7251), .A2(n3350), .B1(n3296), .B2(n1945), .ZN(n5847)
         );
  OAI21_X1 U3935 ( .B1(n4899), .B2(n4900), .A(n3689), .ZN(n4883) );
  OAI221_X1 U3936 ( .B1(n2560), .B2(n3186), .C1(n2552), .C2(n3673), .A(n4902), 
        .ZN(n4899) );
  OAI221_X1 U3937 ( .B1(n2624), .B2(n3226), .C1(n2616), .C2(n3668), .A(n4901), 
        .ZN(n4900) );
  AOI22_X1 U3938 ( .A1(n3168), .A2(n[1025]), .B1(n3153), .B2(n[1033]), .ZN(
        n4902) );
  OAI21_X1 U3939 ( .B1(n4727), .B2(n4728), .A(n3689), .ZN(n4711) );
  OAI221_X1 U3940 ( .B1(n2559), .B2(n3184), .C1(n2551), .C2(n3179), .A(n4730), 
        .ZN(n4727) );
  OAI221_X1 U3941 ( .B1(n2623), .B2(n3218), .C1(n2615), .C2(n3216), .A(n4729), 
        .ZN(n4728) );
  AOI22_X1 U3942 ( .A1(n3168), .A2(n[1026]), .B1(n3154), .B2(n[1034]), .ZN(
        n4730) );
  OAI21_X1 U3943 ( .B1(n4211), .B2(n4212), .A(n3689), .ZN(n4195) );
  OAI221_X1 U3944 ( .B1(n2556), .B2(n3186), .C1(n2548), .C2(n3180), .A(n4214), 
        .ZN(n4211) );
  OAI221_X1 U3945 ( .B1(n2620), .B2(n3221), .C1(n2612), .C2(n3216), .A(n4213), 
        .ZN(n4212) );
  AOI22_X1 U3946 ( .A1(n3164), .A2(n[1029]), .B1(n3156), .B2(n[1037]), .ZN(
        n4214) );
  OAI21_X1 U3947 ( .B1(n4039), .B2(n4040), .A(n3150), .ZN(n4023) );
  OAI221_X1 U3948 ( .B1(n2555), .B2(n3188), .C1(n2547), .C2(n3180), .A(n4042), 
        .ZN(n4039) );
  OAI221_X1 U3949 ( .B1(n2619), .B2(n3223), .C1(n2611), .C2(n3213), .A(n4041), 
        .ZN(n4040) );
  AOI22_X1 U3950 ( .A1(n3166), .A2(n[1030]), .B1(n3155), .B2(n[1038]), .ZN(
        n4042) );
  OAI21_X1 U3951 ( .B1(n4543), .B2(n4544), .A(n3666), .ZN(n4542) );
  OAI221_X1 U3952 ( .B1(n2974), .B2(n3183), .C1(n2966), .C2(n3180), .A(n4546), 
        .ZN(n4543) );
  OAI221_X1 U3953 ( .B1(n3006), .B2(n3667), .C1(n2998), .C2(n3217), .A(n4545), 
        .ZN(n4544) );
  AOI22_X1 U3954 ( .A1(n3164), .A2(n[643]), .B1(n3161), .B2(n[651]), .ZN(n4546) );
  OAI21_X1 U3955 ( .B1(n4563), .B2(n4564), .A(n3698), .ZN(n4562) );
  OAI221_X1 U3956 ( .B1(n3038), .B2(n3187), .C1(n3030), .C2(n3180), .A(n4566), 
        .ZN(n4563) );
  OAI221_X1 U3957 ( .B1(n3070), .B2(n3221), .C1(n3062), .C2(n3217), .A(n4565), 
        .ZN(n4564) );
  AOI22_X1 U3958 ( .A1(n3675), .A2(n[579]), .B1(n3155), .B2(n[587]), .ZN(n4566) );
  OAI21_X1 U3959 ( .B1(n4585), .B2(n4586), .A(n3666), .ZN(n4584) );
  OAI221_X1 U3960 ( .B1(n2302), .B2(n3672), .C1(n2294), .C2(n3180), .A(n4588), 
        .ZN(n4585) );
  OAI221_X1 U3961 ( .B1(n2366), .B2(n3218), .C1(n2358), .C2(n3217), .A(n4587), 
        .ZN(n4586) );
  AOI22_X1 U3962 ( .A1(n3164), .A2(n[1155]), .B1(n3161), .B2(n[1163]), .ZN(
        n4588) );
  OAI21_X1 U3963 ( .B1(n4371), .B2(n4372), .A(n3666), .ZN(n4370) );
  OAI221_X1 U3964 ( .B1(n2973), .B2(n3181), .C1(n2965), .C2(n3673), .A(n4374), 
        .ZN(n4371) );
  OAI221_X1 U3965 ( .B1(n3005), .B2(n3667), .C1(n2997), .C2(n3668), .A(n4373), 
        .ZN(n4372) );
  AOI22_X1 U3966 ( .A1(n3171), .A2(n[644]), .B1(n3676), .B2(n[652]), .ZN(n4374) );
  OAI21_X1 U3967 ( .B1(n4391), .B2(n4392), .A(n3698), .ZN(n4390) );
  OAI221_X1 U3968 ( .B1(n3037), .B2(n3188), .C1(n3029), .C2(n3176), .A(n4394), 
        .ZN(n4391) );
  OAI221_X1 U3969 ( .B1(n3069), .B2(n3226), .C1(n3061), .C2(n3217), .A(n4393), 
        .ZN(n4392) );
  AOI22_X1 U3970 ( .A1(n3163), .A2(n[580]), .B1(n3155), .B2(n[588]), .ZN(n4394) );
  OAI21_X1 U3971 ( .B1(n4413), .B2(n4414), .A(n3666), .ZN(n4412) );
  OAI221_X1 U3972 ( .B1(n2301), .B2(n3672), .C1(n2293), .C2(n3176), .A(n4416), 
        .ZN(n4413) );
  OAI221_X1 U3973 ( .B1(n2365), .B2(n3223), .C1(n2357), .C2(n3217), .A(n4415), 
        .ZN(n4414) );
  AOI22_X1 U3974 ( .A1(n3675), .A2(n[1156]), .B1(n3161), .B2(n[1164]), .ZN(
        n4416) );
  OAI21_X1 U3975 ( .B1(n4433), .B2(n4434), .A(n3698), .ZN(n4432) );
  OAI221_X1 U3976 ( .B1(n2429), .B2(n3184), .C1(n2421), .C2(n3176), .A(n4436), 
        .ZN(n4433) );
  OAI221_X1 U3977 ( .B1(n2493), .B2(n3219), .C1(n2485), .C2(n3213), .A(n4435), 
        .ZN(n4434) );
  AOI22_X1 U3978 ( .A1(n3166), .A2(n[1092]), .B1(n3161), .B2(n[1100]), .ZN(
        n4436) );
  OAI21_X1 U3979 ( .B1(n4455), .B2(n4456), .A(n3666), .ZN(n4454) );
  OAI221_X1 U3980 ( .B1(n1277), .B2(n3189), .C1(n1269), .C2(n3173), .A(n4458), 
        .ZN(n4455) );
  OAI221_X1 U3981 ( .B1(n1341), .B2(n3225), .C1(n1333), .C2(n3211), .A(n4457), 
        .ZN(n4456) );
  AOI22_X1 U3982 ( .A1(n3165), .A2(n[1668]), .B1(n3161), .B2(n[1676]), .ZN(
        n4458) );
  OAI21_X1 U3983 ( .B1(n4475), .B2(n4476), .A(n3698), .ZN(n4474) );
  OAI221_X1 U3984 ( .B1(n1405), .B2(n3186), .C1(n1397), .C2(n3180), .A(n4478), 
        .ZN(n4475) );
  OAI221_X1 U3985 ( .B1(n1469), .B2(n3226), .C1(n1461), .C2(n3215), .A(n4477), 
        .ZN(n4476) );
  AOI22_X1 U3986 ( .A1(n3171), .A2(n[1604]), .B1(n3154), .B2(n[1612]), .ZN(
        n4478) );
  OAI21_X1 U3987 ( .B1(n4497), .B2(n4498), .A(n3666), .ZN(n4496) );
  OAI221_X1 U3988 ( .B1(n413), .B2(n3672), .C1(n405), .C2(n3175), .A(n4500), 
        .ZN(n4497) );
  OAI221_X1 U3989 ( .B1(n445), .B2(n3667), .C1(n437), .C2(n3214), .A(n4499), 
        .ZN(n4498) );
  AOI22_X1 U3990 ( .A1(n3171), .A2(n[2180]), .B1(n3159), .B2(n[2188]), .ZN(
        n4500) );
  OAI21_X1 U3991 ( .B1(n4517), .B2(n4518), .A(n3698), .ZN(n4516) );
  OAI221_X1 U3992 ( .B1(n477), .B2(n3189), .C1(n469), .C2(n3180), .A(n4520), 
        .ZN(n4517) );
  OAI221_X1 U3993 ( .B1(n509), .B2(n3220), .C1(n501), .C2(n3217), .A(n4519), 
        .ZN(n4518) );
  AOI22_X1 U3994 ( .A1(n3171), .A2(n[2116]), .B1(n3154), .B2(n[2124]), .ZN(
        n4520) );
  OAI21_X1 U3995 ( .B1(n4345), .B2(n4346), .A(n3698), .ZN(n4344) );
  OAI221_X1 U3996 ( .B1(n476), .B2(n3185), .C1(n468), .C2(n3176), .A(n4348), 
        .ZN(n4345) );
  OAI221_X1 U3997 ( .B1(n508), .B2(n3218), .C1(n500), .C2(n3214), .A(n4347), 
        .ZN(n4346) );
  AOI22_X1 U3998 ( .A1(n3170), .A2(n[2117]), .B1(n3160), .B2(n[2125]), .ZN(
        n4348) );
  OAI21_X1 U3999 ( .B1(n3897), .B2(n3898), .A(n3666), .ZN(n3896) );
  OAI221_X1 U4000 ( .B1(n2298), .B2(n3672), .C1(n2290), .C2(n3176), .A(n3900), 
        .ZN(n3897) );
  OAI221_X1 U4001 ( .B1(n2362), .B2(n3218), .C1(n2354), .C2(n3213), .A(n3899), 
        .ZN(n3898) );
  AOI22_X1 U4002 ( .A1(n3162), .A2(n[1159]), .B1(n3157), .B2(n[1167]), .ZN(
        n3900) );
  OAI21_X1 U4003 ( .B1(n3917), .B2(n3918), .A(n3698), .ZN(n3916) );
  OAI221_X1 U4004 ( .B1(n2426), .B2(n3181), .C1(n2418), .C2(n3176), .A(n3920), 
        .ZN(n3917) );
  OAI221_X1 U4005 ( .B1(n2490), .B2(n3219), .C1(n2482), .C2(n3213), .A(n3919), 
        .ZN(n3918) );
  AOI22_X1 U4006 ( .A1(n3169), .A2(n[1095]), .B1(n3157), .B2(n[1103]), .ZN(
        n3920) );
  OAI21_X1 U4007 ( .B1(n3939), .B2(n3940), .A(n3666), .ZN(n3938) );
  OAI221_X1 U4008 ( .B1(n1274), .B2(n3181), .C1(n1266), .C2(n3176), .A(n3942), 
        .ZN(n3939) );
  OAI221_X1 U4009 ( .B1(n1338), .B2(n3221), .C1(n1330), .C2(n3213), .A(n3941), 
        .ZN(n3940) );
  AOI22_X1 U4010 ( .A1(n3162), .A2(n[1671]), .B1(n3157), .B2(n[1679]), .ZN(
        n3942) );
  OAI21_X1 U4011 ( .B1(n3855), .B2(n3856), .A(n3227), .ZN(n3854) );
  OAI221_X1 U4012 ( .B1(n2970), .B2(n3672), .C1(n2962), .C2(n3177), .A(n3858), 
        .ZN(n3855) );
  OAI221_X1 U4013 ( .B1(n3002), .B2(n3225), .C1(n2994), .C2(n3214), .A(n3857), 
        .ZN(n3856) );
  AOI22_X1 U4014 ( .A1(n3168), .A2(n[647]), .B1(n3158), .B2(n[655]), .ZN(n3858) );
  OAI21_X1 U4015 ( .B1(n3875), .B2(n3876), .A(n3149), .ZN(n3874) );
  OAI221_X1 U4016 ( .B1(n3034), .B2(n3185), .C1(n3026), .C2(n3177), .A(n3878), 
        .ZN(n3875) );
  OAI221_X1 U4017 ( .B1(n3066), .B2(n3225), .C1(n3058), .C2(n3214), .A(n3877), 
        .ZN(n3876) );
  AOI22_X1 U4018 ( .A1(n3168), .A2(n[583]), .B1(n3158), .B2(n[591]), .ZN(n3878) );
  OAI21_X1 U4019 ( .B1(n3723), .B2(n3724), .A(n3666), .ZN(n3722) );
  OAI221_X1 U4020 ( .B1(n2297), .B2(n3184), .C1(n2289), .C2(n3179), .A(n3726), 
        .ZN(n3723) );
  OAI221_X1 U4021 ( .B1(n2361), .B2(n3222), .C1(n2353), .C2(n3216), .A(n3725), 
        .ZN(n3724) );
  AOI22_X1 U4022 ( .A1(n3170), .A2(n[1160]), .B1(n3160), .B2(n[1168]), .ZN(
        n3726) );
  OAI21_X1 U4023 ( .B1(n3743), .B2(n3744), .A(n3698), .ZN(n3742) );
  OAI221_X1 U4024 ( .B1(n2425), .B2(n3181), .C1(n2417), .C2(n3179), .A(n3746), 
        .ZN(n3743) );
  OAI221_X1 U4025 ( .B1(n2489), .B2(n3226), .C1(n2481), .C2(n3216), .A(n3745), 
        .ZN(n3744) );
  AOI22_X1 U4026 ( .A1(n3170), .A2(n[1096]), .B1(n3160), .B2(n[1104]), .ZN(
        n3746) );
  OAI21_X1 U4027 ( .B1(n3766), .B2(n3767), .A(n3666), .ZN(n3765) );
  OAI221_X1 U4028 ( .B1(n1273), .B2(n3182), .C1(n1265), .C2(n3178), .A(n3769), 
        .ZN(n3766) );
  OAI221_X1 U4029 ( .B1(n1337), .B2(n3222), .C1(n1329), .C2(n3215), .A(n3768), 
        .ZN(n3767) );
  AOI22_X1 U4030 ( .A1(n3169), .A2(n[1672]), .B1(n3159), .B2(n[1680]), .ZN(
        n3769) );
  OAI21_X1 U4031 ( .B1(n3786), .B2(n3787), .A(n3698), .ZN(n3785) );
  OAI221_X1 U4032 ( .B1(n1401), .B2(n3183), .C1(n1393), .C2(n3178), .A(n3789), 
        .ZN(n3786) );
  OAI221_X1 U4033 ( .B1(n1465), .B2(n3220), .C1(n1457), .C2(n3215), .A(n3788), 
        .ZN(n3787) );
  AOI22_X1 U4034 ( .A1(n3169), .A2(n[1608]), .B1(n3159), .B2(n[1616]), .ZN(
        n3789) );
  OAI21_X1 U4035 ( .B1(n3696), .B2(n3697), .A(n3149), .ZN(n3695) );
  OAI221_X1 U4036 ( .B1(n3033), .B2(n3672), .C1(n3025), .C2(n3179), .A(n3700), 
        .ZN(n3696) );
  OAI221_X1 U4037 ( .B1(n3065), .B2(n3224), .C1(n3057), .C2(n3216), .A(n3699), 
        .ZN(n3697) );
  AOI22_X1 U4038 ( .A1(n3170), .A2(n[584]), .B1(n3160), .B2(n[592]), .ZN(n3700) );
  OAI21_X1 U4039 ( .B1(n3664), .B2(n3665), .A(n3227), .ZN(n3663) );
  OAI221_X1 U4040 ( .B1(n2969), .B2(n3188), .C1(n2961), .C2(n3180), .A(n3674), 
        .ZN(n3664) );
  OAI221_X1 U4041 ( .B1(n3001), .B2(n3226), .C1(n2993), .C2(n3217), .A(n3669), 
        .ZN(n3665) );
  AOI22_X1 U4042 ( .A1(n3171), .A2(n[648]), .B1(n3161), .B2(n[656]), .ZN(n3674) );
  OAI21_X1 U4043 ( .B1(n3809), .B2(n3810), .A(n3666), .ZN(n3808) );
  OAI221_X1 U4044 ( .B1(n409), .B2(n3184), .C1(n401), .C2(n3178), .A(n3812), 
        .ZN(n3809) );
  OAI221_X1 U4045 ( .B1(n441), .B2(n3218), .C1(n433), .C2(n3215), .A(n3811), 
        .ZN(n3810) );
  AOI22_X1 U4046 ( .A1(n3169), .A2(n[2184]), .B1(n3159), .B2(n[2192]), .ZN(
        n3812) );
  OAI21_X1 U4047 ( .B1(n3829), .B2(n3830), .A(n3698), .ZN(n3828) );
  OAI221_X1 U4048 ( .B1(n473), .B2(n3183), .C1(n465), .C2(n3177), .A(n3832), 
        .ZN(n3829) );
  OAI221_X1 U4049 ( .B1(n505), .B2(n3225), .C1(n497), .C2(n3214), .A(n3831), 
        .ZN(n3830) );
  AOI22_X1 U4050 ( .A1(n3168), .A2(n[2120]), .B1(n3158), .B2(n[2128]), .ZN(
        n3832) );
  OAI21_X1 U4051 ( .B1(n4547), .B2(n4548), .A(n3679), .ZN(n4541) );
  OAI221_X1 U4052 ( .B1(n2846), .B2(n3182), .C1(n2838), .C2(n3180), .A(n4550), 
        .ZN(n4547) );
  OAI221_X1 U4053 ( .B1(n2878), .B2(n3225), .C1(n2870), .C2(n3217), .A(n4549), 
        .ZN(n4548) );
  AOI22_X1 U4054 ( .A1(n3675), .A2(n[771]), .B1(n3153), .B2(n[779]), .ZN(n4550) );
  OAI21_X1 U4055 ( .B1(n4567), .B2(n4568), .A(n3148), .ZN(n4561) );
  OAI221_X1 U4056 ( .B1(n2910), .B2(n3186), .C1(n2902), .C2(n3173), .A(n4570), 
        .ZN(n4567) );
  OAI221_X1 U4057 ( .B1(n2942), .B2(n3223), .C1(n2934), .C2(n3216), .A(n4569), 
        .ZN(n4568) );
  AOI22_X1 U4058 ( .A1(n3165), .A2(n[707]), .B1(n3160), .B2(n[715]), .ZN(n4570) );
  OAI21_X1 U4059 ( .B1(n4375), .B2(n4376), .A(n3679), .ZN(n4369) );
  OAI221_X1 U4060 ( .B1(n2845), .B2(n3181), .C1(n2837), .C2(n3172), .A(n4378), 
        .ZN(n4375) );
  OAI221_X1 U4061 ( .B1(n2877), .B2(n3667), .C1(n2869), .C2(n3209), .A(n4377), 
        .ZN(n4376) );
  AOI22_X1 U4062 ( .A1(n3164), .A2(n[772]), .B1(n3153), .B2(n[780]), .ZN(n4378) );
  OAI21_X1 U4063 ( .B1(n4395), .B2(n4396), .A(n3148), .ZN(n4389) );
  OAI221_X1 U4064 ( .B1(n2909), .B2(n3672), .C1(n2901), .C2(n3175), .A(n4398), 
        .ZN(n4395) );
  OAI221_X1 U4065 ( .B1(n2941), .B2(n3222), .C1(n2933), .C2(n3668), .A(n4397), 
        .ZN(n4396) );
  AOI22_X1 U4066 ( .A1(n3171), .A2(n[708]), .B1(n3160), .B2(n[716]), .ZN(n4398) );
  OAI21_X1 U4067 ( .B1(n3901), .B2(n3902), .A(n3679), .ZN(n3895) );
  OAI221_X1 U4068 ( .B1(n2042), .B2(n3181), .C1(n2034), .C2(n3176), .A(n3904), 
        .ZN(n3901) );
  OAI221_X1 U4069 ( .B1(n2106), .B2(n3224), .C1(n2098), .C2(n3213), .A(n3903), 
        .ZN(n3902) );
  AOI22_X1 U4070 ( .A1(n3171), .A2(n[1287]), .B1(n3157), .B2(n[1295]), .ZN(
        n3904) );
  OAI21_X1 U4071 ( .B1(n3921), .B2(n3922), .A(n3703), .ZN(n3915) );
  OAI221_X1 U4072 ( .B1(n2170), .B2(n3181), .C1(n2162), .C2(n3176), .A(n3924), 
        .ZN(n3921) );
  OAI221_X1 U4073 ( .B1(n2234), .B2(n3224), .C1(n2226), .C2(n3213), .A(n3923), 
        .ZN(n3922) );
  AOI22_X1 U4074 ( .A1(n3166), .A2(n[1223]), .B1(n3157), .B2(n[1231]), .ZN(
        n3924) );
  OAI21_X1 U4075 ( .B1(n3727), .B2(n3728), .A(n3679), .ZN(n3721) );
  OAI221_X1 U4076 ( .B1(n2041), .B2(n3188), .C1(n2033), .C2(n3179), .A(n3730), 
        .ZN(n3727) );
  OAI221_X1 U4077 ( .B1(n2105), .B2(n3221), .C1(n2097), .C2(n3216), .A(n3729), 
        .ZN(n3728) );
  AOI22_X1 U4078 ( .A1(n3170), .A2(n[1288]), .B1(n3160), .B2(n[1296]), .ZN(
        n3730) );
  OAI21_X1 U4079 ( .B1(n3747), .B2(n3748), .A(n3703), .ZN(n3741) );
  OAI221_X1 U4080 ( .B1(n2169), .B2(n3672), .C1(n2161), .C2(n3179), .A(n3750), 
        .ZN(n3747) );
  OAI221_X1 U4081 ( .B1(n2233), .B2(n3220), .C1(n2225), .C2(n3216), .A(n3749), 
        .ZN(n3748) );
  AOI22_X1 U4082 ( .A1(n3170), .A2(n[1224]), .B1(n3160), .B2(n[1232]), .ZN(
        n3750) );
  OAI21_X1 U4083 ( .B1(n4551), .B2(n4552), .A(n3684), .ZN(n4540) );
  OAI221_X1 U4084 ( .B1(n2718), .B2(n3185), .C1(n2710), .C2(n3180), .A(n4554), 
        .ZN(n4551) );
  OAI221_X1 U4085 ( .B1(n2750), .B2(n3221), .C1(n2742), .C2(n3217), .A(n4553), 
        .ZN(n4552) );
  AOI22_X1 U4086 ( .A1(n3170), .A2(n[899]), .B1(n3160), .B2(n[907]), .ZN(n4554) );
  OAI21_X1 U4087 ( .B1(n4571), .B2(n4572), .A(n3708), .ZN(n4560) );
  OAI221_X1 U4088 ( .B1(n2782), .B2(n3188), .C1(n2774), .C2(n3176), .A(n4574), 
        .ZN(n4571) );
  OAI221_X1 U4089 ( .B1(n2814), .B2(n3219), .C1(n2806), .C2(n3213), .A(n4573), 
        .ZN(n4572) );
  AOI22_X1 U4090 ( .A1(n3165), .A2(n[835]), .B1(n3676), .B2(n[843]), .ZN(n4574) );
  OAI21_X1 U4091 ( .B1(n4379), .B2(n4380), .A(n3684), .ZN(n4368) );
  OAI221_X1 U4092 ( .B1(n2717), .B2(n3183), .C1(n2709), .C2(n3673), .A(n4382), 
        .ZN(n4379) );
  OAI221_X1 U4093 ( .B1(n2749), .B2(n3224), .C1(n2741), .C2(n3668), .A(n4381), 
        .ZN(n4380) );
  AOI22_X1 U4094 ( .A1(n3170), .A2(n[900]), .B1(n3161), .B2(n[908]), .ZN(n4382) );
  OAI21_X1 U4095 ( .B1(n4399), .B2(n4400), .A(n3708), .ZN(n4388) );
  OAI221_X1 U4096 ( .B1(n2781), .B2(n3182), .C1(n2773), .C2(n3673), .A(n4402), 
        .ZN(n4399) );
  OAI221_X1 U4097 ( .B1(n2813), .B2(n3219), .C1(n2805), .C2(n3211), .A(n4401), 
        .ZN(n4400) );
  AOI22_X1 U4098 ( .A1(n3164), .A2(n[836]), .B1(n3157), .B2(n[844]), .ZN(n4402) );
  OAI21_X1 U4099 ( .B1(n3905), .B2(n3906), .A(n3684), .ZN(n3894) );
  OAI221_X1 U4100 ( .B1(n1786), .B2(n3181), .C1(n1778), .C2(n3176), .A(n3908), 
        .ZN(n3905) );
  OAI221_X1 U4101 ( .B1(n1850), .B2(n3219), .C1(n1842), .C2(n3213), .A(n3907), 
        .ZN(n3906) );
  AOI22_X1 U4102 ( .A1(n3163), .A2(n[1415]), .B1(n3157), .B2(n[1423]), .ZN(
        n3908) );
  OAI21_X1 U4103 ( .B1(n3925), .B2(n3926), .A(n3708), .ZN(n3914) );
  OAI221_X1 U4104 ( .B1(n1914), .B2(n3181), .C1(n1906), .C2(n3176), .A(n3928), 
        .ZN(n3925) );
  OAI221_X1 U4105 ( .B1(n1978), .B2(n3218), .C1(n1970), .C2(n3213), .A(n3927), 
        .ZN(n3926) );
  AOI22_X1 U4106 ( .A1(n3162), .A2(n[1351]), .B1(n3157), .B2(n[1359]), .ZN(
        n3928) );
  OAI21_X1 U4107 ( .B1(n3731), .B2(n3732), .A(n3684), .ZN(n3720) );
  OAI221_X1 U4108 ( .B1(n1785), .B2(n3181), .C1(n1777), .C2(n3179), .A(n3734), 
        .ZN(n3731) );
  OAI221_X1 U4109 ( .B1(n1849), .B2(n3218), .C1(n1841), .C2(n3216), .A(n3733), 
        .ZN(n3732) );
  AOI22_X1 U4110 ( .A1(n3170), .A2(n[1416]), .B1(n3160), .B2(n[1424]), .ZN(
        n3734) );
  OAI21_X1 U4111 ( .B1(n3751), .B2(n3752), .A(n3708), .ZN(n3740) );
  OAI221_X1 U4112 ( .B1(n1913), .B2(n3672), .C1(n1905), .C2(n3179), .A(n3754), 
        .ZN(n3751) );
  OAI221_X1 U4113 ( .B1(n1977), .B2(n3218), .C1(n1969), .C2(n3216), .A(n3753), 
        .ZN(n3752) );
  AOI22_X1 U4114 ( .A1(n3170), .A2(n[1352]), .B1(n3160), .B2(n[1360]), .ZN(
        n3754) );
  OAI21_X1 U4115 ( .B1(n4555), .B2(n4556), .A(n3689), .ZN(n4539) );
  OAI221_X1 U4116 ( .B1(n2558), .B2(n3672), .C1(n2550), .C2(n3175), .A(n4558), 
        .ZN(n4555) );
  OAI221_X1 U4117 ( .B1(n2622), .B2(n3218), .C1(n2614), .C2(n3217), .A(n4557), 
        .ZN(n4556) );
  AOI22_X1 U4118 ( .A1(n3162), .A2(n[1027]), .B1(n3676), .B2(n[1035]), .ZN(
        n4558) );
  OAI21_X1 U4119 ( .B1(n4383), .B2(n4384), .A(n3689), .ZN(n4367) );
  OAI221_X1 U4120 ( .B1(n2557), .B2(n3189), .C1(n2549), .C2(n3174), .A(n4386), 
        .ZN(n4383) );
  OAI221_X1 U4121 ( .B1(n2621), .B2(n3225), .C1(n2613), .C2(n3217), .A(n4385), 
        .ZN(n4384) );
  AOI22_X1 U4122 ( .A1(n3165), .A2(n[1028]), .B1(n3158), .B2(n[1036]), .ZN(
        n4386) );
  OAI21_X1 U4123 ( .B1(n3909), .B2(n3910), .A(n3150), .ZN(n3893) );
  OAI221_X1 U4124 ( .B1(n1530), .B2(n3181), .C1(n1522), .C2(n3176), .A(n3912), 
        .ZN(n3909) );
  OAI221_X1 U4125 ( .B1(n1594), .B2(n3225), .C1(n1586), .C2(n3213), .A(n3911), 
        .ZN(n3910) );
  AOI22_X1 U4126 ( .A1(n3163), .A2(n[1543]), .B1(n3157), .B2(n[1551]), .ZN(
        n3912) );
  OAI21_X1 U4127 ( .B1(n3735), .B2(n3736), .A(n3150), .ZN(n3719) );
  OAI221_X1 U4128 ( .B1(n1529), .B2(n3672), .C1(n1521), .C2(n3179), .A(n3738), 
        .ZN(n3735) );
  OAI221_X1 U4129 ( .B1(n1593), .B2(n3219), .C1(n1585), .C2(n3216), .A(n3737), 
        .ZN(n3736) );
  AOI22_X1 U4130 ( .A1(n3170), .A2(n[1544]), .B1(n3160), .B2(n[1552]), .ZN(
        n3738) );
  INV_X1 U4131 ( .A(data_w[0]), .ZN(n7258) );
  INV_X1 U4132 ( .A(data_w[1]), .ZN(n7257) );
  INV_X1 U4133 ( .A(data_w[2]), .ZN(n7256) );
  INV_X1 U4134 ( .A(data_w[3]), .ZN(n7255) );
  INV_X1 U4135 ( .A(data_w[4]), .ZN(n7254) );
  INV_X1 U4136 ( .A(data_w[5]), .ZN(n7253) );
  INV_X1 U4137 ( .A(data_w[6]), .ZN(n7252) );
  INV_X1 U4138 ( .A(data_w[7]), .ZN(n7251) );
  BUF_X1 U4139 ( .A(n7251), .Z(n3074) );
  BUF_X1 U4140 ( .A(n7252), .Z(n3083) );
  BUF_X1 U4141 ( .A(n7253), .Z(n3092) );
  BUF_X1 U4142 ( .A(n7256), .Z(n3119) );
  BUF_X1 U4143 ( .A(n7257), .Z(n3130) );
  BUF_X1 U4144 ( .A(n7258), .Z(n3138) );
  BUF_X1 U4145 ( .A(n3153), .Z(n3154) );
  BUF_X1 U4146 ( .A(n3153), .Z(n3155) );
  BUF_X1 U4147 ( .A(n3153), .Z(n3156) );
  BUF_X1 U4148 ( .A(n3153), .Z(n3157) );
  BUF_X1 U4149 ( .A(n3153), .Z(n3161) );
  BUF_X1 U4150 ( .A(n3675), .Z(n3162) );
  BUF_X1 U4151 ( .A(n3675), .Z(n3163) );
  BUF_X1 U4152 ( .A(n3675), .Z(n3164) );
  BUF_X1 U4153 ( .A(n3675), .Z(n3165) );
  BUF_X1 U4154 ( .A(n3675), .Z(n3166) );
  BUF_X1 U4155 ( .A(n3675), .Z(n3167) );
  BUF_X1 U4156 ( .A(n3675), .Z(n3171) );
  BUF_X1 U4157 ( .A(n3172), .Z(n3173) );
  BUF_X1 U4158 ( .A(n3172), .Z(n3174) );
  BUF_X1 U4159 ( .A(n3172), .Z(n3175) );
  BUF_X1 U4160 ( .A(n3172), .Z(n3180) );
  BUF_X1 U4161 ( .A(n3672), .Z(n3182) );
  BUF_X1 U4162 ( .A(n3672), .Z(n3183) );
  BUF_X1 U4163 ( .A(n3181), .Z(n3184) );
  BUF_X1 U4164 ( .A(n3181), .Z(n3185) );
  BUF_X1 U4165 ( .A(n3181), .Z(n3186) );
  BUF_X1 U4166 ( .A(n3181), .Z(n3187) );
  BUF_X1 U4167 ( .A(n3181), .Z(n3188) );
  BUF_X1 U4168 ( .A(n3181), .Z(n3189) );
  BUF_X1 U4169 ( .A(n3671), .Z(n3191) );
  BUF_X1 U4170 ( .A(n3671), .Z(n3192) );
  BUF_X1 U4171 ( .A(n3190), .Z(n3193) );
  BUF_X1 U4172 ( .A(n3190), .Z(n3194) );
  BUF_X1 U4173 ( .A(n3190), .Z(n3195) );
  BUF_X1 U4174 ( .A(n3190), .Z(n3196) );
  BUF_X1 U4175 ( .A(n3190), .Z(n3197) );
  BUF_X1 U4176 ( .A(n3190), .Z(n3198) );
  BUF_X1 U4177 ( .A(n3670), .Z(n3199) );
  BUF_X1 U4178 ( .A(n3670), .Z(n3200) );
  BUF_X1 U4179 ( .A(n3670), .Z(n3201) );
  BUF_X1 U4180 ( .A(n3670), .Z(n3202) );
  BUF_X1 U4181 ( .A(n3670), .Z(n3203) );
  BUF_X1 U4182 ( .A(n3670), .Z(n3204) );
  BUF_X1 U4183 ( .A(n3670), .Z(n3208) );
  BUF_X1 U4184 ( .A(n3209), .Z(n3210) );
  BUF_X1 U4185 ( .A(n3209), .Z(n3211) );
  BUF_X1 U4186 ( .A(n3209), .Z(n3212) );
  BUF_X1 U4187 ( .A(n3209), .Z(n3217) );
  BUF_X1 U4188 ( .A(n3667), .Z(n3218) );
  BUF_X1 U4189 ( .A(n3667), .Z(n3219) );
  BUF_X1 U4190 ( .A(n3667), .Z(n3220) );
  BUF_X1 U4191 ( .A(n3667), .Z(n3221) );
  BUF_X1 U4192 ( .A(n3667), .Z(n3222) );
  BUF_X1 U4193 ( .A(n3667), .Z(n3223) );
  BUF_X1 U4194 ( .A(n3667), .Z(n3224) );
  BUF_X1 U4195 ( .A(n3667), .Z(n3226) );
endmodule


module asyn_fifo_top_word_width8_0 ( r_clk, w_clk, rd, wr, reset_n, data_in, 
        data_out, full, empty );
  input [7:0] data_in;
  output [7:0] data_out;
  input r_clk, w_clk, rd, wr, reset_n;
  output full, empty;
  wire   we_enable;
  wire   [7:0] addr_r;
  wire   [7:0] addr_w;

  fifo_control_unit_addr_size8_0 fifo_ctrl ( .reset_n(reset_n), .w_clk(w_clk), 
        .r_clk(r_clk), .rd(rd), .wr(wr), .addr_r(addr_r), .addr_w(addr_w), 
        .full(full), .empty(empty), .we_enable(we_enable) );
  reg_memory_file_addr_size8_word_width8_0 fifo_memory ( .we_s(we_enable), 
        .clk(w_clk), .addr_r(addr_r), .addr_w(addr_w), .data_w(data_in), 
        .data_r(data_out) );
endmodule


module timer_bits10 ( clk, enable, reset, final, tkl );
  input [9:0] final;
  input clk, enable, reset;
  output tkl;
  wire   n1, n2, n3, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n19,
         n21, n22, n23, n24, n25, n26, n29, n31, n32, n35, n36, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n67, n68, n69,
         n70, n71, n72, n66, n73, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84;

  XOR2_X1 U4 ( .A(n60), .B(n3), .Z(n2) );
  XOR2_X1 U56 ( .A(n51), .B(final[4]), .Z(n46) );
  DFFR_X1 Q_reg_reg_10_ ( .D(n62), .CK(clk), .RN(reset), .QN(n60) );
  DFFR_X1 Q_reg_reg_9_ ( .D(n63), .CK(clk), .RN(reset), .QN(n59) );
  DFFR_X1 Q_reg_reg_8_ ( .D(n64), .CK(clk), .RN(reset), .QN(n58) );
  DFFR_X1 Q_reg_reg_5_ ( .D(n67), .CK(clk), .RN(reset), .Q(n82), .QN(n56) );
  DFFR_X1 Q_reg_reg_1_ ( .D(n71), .CK(clk), .RN(reset), .QN(n54) );
  DFFR_X1 Q_reg_reg_0_ ( .D(n72), .CK(clk), .RN(reset), .Q(n77), .QN(n61) );
  DFFR_X1 Q_reg_reg_2_ ( .D(n70), .CK(clk), .RN(reset), .Q(n80), .QN(n53) );
  DFFR_X1 Q_reg_reg_6_ ( .D(n73), .CK(clk), .RN(reset), .Q(n83), .QN(n55) );
  DFFR_X1 Q_reg_reg_7_ ( .D(n65), .CK(clk), .RN(reset), .QN(n57) );
  DFFR_X1 Q_reg_reg_3_ ( .D(n69), .CK(clk), .RN(reset), .Q(n81), .QN(n52) );
  DFFR_X1 Q_reg_reg_4_ ( .D(n68), .CK(clk), .RN(reset), .QN(n51) );
  INV_X1 U3 ( .A(n9), .ZN(tkl) );
  AOI21_X1 U5 ( .B1(n9), .B2(n78), .A(n84), .ZN(n21) );
  OAI21_X1 U6 ( .B1(tkl), .B2(n80), .A(n32), .ZN(n29) );
  NOR2_X1 U7 ( .A1(n84), .A2(n9), .ZN(n1) );
  INV_X1 U8 ( .A(n10), .ZN(n78) );
  INV_X1 U9 ( .A(n6), .ZN(n79) );
  NAND4_X1 U10 ( .A1(n60), .A2(n38), .A3(n39), .A4(n40), .ZN(n9) );
  XNOR2_X1 U11 ( .A(n77), .B(final[0]), .ZN(n38) );
  NOR3_X1 U12 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n39) );
  NOR4_X1 U13 ( .A1(n41), .A2(n42), .A3(n43), .A4(n44), .ZN(n40) );
  XNOR2_X1 U14 ( .A(n54), .B(final[1]), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n56), .B(final[5]), .ZN(n49) );
  XNOR2_X1 U16 ( .A(n55), .B(final[6]), .ZN(n43) );
  XNOR2_X1 U17 ( .A(n57), .B(final[7]), .ZN(n50) );
  XNOR2_X1 U18 ( .A(n58), .B(final[8]), .ZN(n42) );
  NAND3_X1 U19 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n41) );
  XNOR2_X1 U20 ( .A(n81), .B(final[3]), .ZN(n45) );
  XNOR2_X1 U21 ( .A(n80), .B(final[2]), .ZN(n47) );
  XNOR2_X1 U22 ( .A(n59), .B(final[9]), .ZN(n48) );
  NOR3_X1 U23 ( .A1(n61), .A2(n54), .A3(n19), .ZN(n26) );
  NOR3_X1 U24 ( .A1(n78), .A2(n56), .A3(n19), .ZN(n15) );
  AOI21_X1 U25 ( .B1(n9), .B2(n61), .A(n84), .ZN(n35) );
  AOI21_X1 U26 ( .B1(n9), .B2(n54), .A(n76), .ZN(n32) );
  INV_X1 U27 ( .A(n35), .ZN(n76) );
  NAND2_X1 U28 ( .A1(enable), .A2(n9), .ZN(n19) );
  OAI21_X1 U29 ( .B1(tkl), .B2(n82), .A(n21), .ZN(n16) );
  OAI22_X1 U30 ( .A1(n53), .A2(n32), .B1(n80), .B2(n75), .ZN(n70) );
  INV_X1 U31 ( .A(n26), .ZN(n75) );
  OAI21_X1 U32 ( .B1(n52), .B2(n66), .A(n31), .ZN(n69) );
  NAND3_X1 U33 ( .A1(n52), .A2(n80), .A3(n26), .ZN(n31) );
  INV_X1 U34 ( .A(n29), .ZN(n66) );
  OAI21_X1 U35 ( .B1(n57), .B2(n12), .A(n13), .ZN(n65) );
  NAND3_X1 U36 ( .A1(n57), .A2(n83), .A3(n15), .ZN(n13) );
  AOI21_X1 U37 ( .B1(n55), .B2(n9), .A(n16), .ZN(n12) );
  OAI21_X1 U38 ( .B1(n51), .B2(n24), .A(n25), .ZN(n68) );
  NAND4_X1 U39 ( .A1(n26), .A2(n51), .A3(n80), .A4(n81), .ZN(n25) );
  AOI21_X1 U40 ( .B1(n52), .B2(n9), .A(n29), .ZN(n24) );
  INV_X1 U41 ( .A(n17), .ZN(n73) );
  AOI22_X1 U42 ( .A1(n83), .A2(n16), .B1(n55), .B2(n15), .ZN(n17) );
  AOI211_X1 U43 ( .C1(n58), .C2(n7), .A(n1), .B(n6), .ZN(n64) );
  OAI22_X1 U44 ( .A1(n56), .A2(n21), .B1(n19), .B2(n22), .ZN(n67) );
  NAND2_X1 U45 ( .A1(n10), .A2(n56), .ZN(n22) );
  OAI22_X1 U46 ( .A1(n54), .A2(n35), .B1(n19), .B2(n36), .ZN(n71) );
  NAND2_X1 U47 ( .A1(n54), .A2(n77), .ZN(n36) );
  OAI22_X1 U48 ( .A1(n61), .A2(enable), .B1(n77), .B2(n19), .ZN(n72) );
  NOR2_X1 U49 ( .A1(n1), .A2(n2), .ZN(n62) );
  NOR2_X1 U50 ( .A1(n59), .A2(n79), .ZN(n3) );
  NOR2_X1 U51 ( .A1(n1), .A2(n5), .ZN(n63) );
  XNOR2_X1 U52 ( .A(n59), .B(n79), .ZN(n5) );
  NOR4_X1 U53 ( .A1(n61), .A2(n54), .A3(n23), .A4(n53), .ZN(n10) );
  OR2_X1 U54 ( .A1(n51), .A2(n52), .ZN(n23) );
  NAND3_X1 U55 ( .A1(n10), .A2(enable), .A3(n11), .ZN(n7) );
  NOR3_X1 U57 ( .A1(n57), .A2(n55), .A3(n56), .ZN(n11) );
  NOR2_X1 U58 ( .A1(n7), .A2(n58), .ZN(n6) );
  INV_X1 U59 ( .A(enable), .ZN(n84) );
endmodule


module UART ( clk, reset_n, wr_uart, data_w, tx, tx_full, rx, rd_uart, data_r, 
        rx_empty, rx_err, rx_done, fr_err, baud_final );
  input [7:0] data_w;
  output [7:0] data_r;
  input [9:0] baud_final;
  input clk, reset_n, wr_uart, rx, rd_uart;
  output tx, tx_full, rx_empty, rx_err, rx_done, fr_err;
  wire   s_tick, tx_done, empty, n2;
  wire   [7:0] data_in;
  wire   [7:0] data_out;

  tx_D_bits9_sb_tick16 Uart_transmitter ( .clk(clk), .reset_n(reset_n), 
        .data_in(data_in), .tx_start(n2), .s_tick(s_tick), .tx(tx), .tx_done(
        tx_done) );
  asyn_fifo_top_word_width8_1 tx_fifo ( .r_clk(clk), .w_clk(clk), .rd(tx_done), 
        .wr(wr_uart), .reset_n(reset_n), .data_in(data_w), .data_out(data_in), 
        .full(tx_full), .empty(empty) );
  rx_D_bits9_sb_tick16 Uart_reciever ( .clk(clk), .reset_n(reset_n), .rx(rx), 
        .s_tick(s_tick), .data_out(data_out), .rx_done(rx_done), .rx_err(
        rx_err), .fr_err(fr_err) );
  asyn_fifo_top_word_width8_0 rx_fifo ( .r_clk(clk), .w_clk(clk), .rd(rd_uart), 
        .wr(rx_done), .reset_n(reset_n), .data_in(data_out), .data_out(data_r), 
        .empty(rx_empty) );
  timer_bits10 baud_rate ( .clk(clk), .enable(1'b1), .reset(reset_n), .final(
        baud_final), .tkl(s_tick) );
  INV_X1 U3 ( .A(empty), .ZN(n2) );
endmodule

